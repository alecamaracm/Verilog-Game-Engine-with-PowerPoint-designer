module PP2VerilogDrawingController(xPixel,yPixel,VGAr,VGAg,VGAb);

input [9:0]xPixel;
input[8:0]yPixel;
output [7:0]VGAr;
output [7:0]VGAg;
output [7:0]VGAb;
reg [7:0]VGAr;
reg [7:0]VGAg;
reg [7:0]VGAb;

always @(*)
begin

	//Writing backgound color
	VGAr = 8'b11111111;
	VGAg = 8'b11111111; 
	VGAb = 8'b11111111; 

	//Drawing picture with compression rate: 1:1
	if(xPixel>=0 && xPixel<1 && yPixel>=0 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=124 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=147 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=253 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=271 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=278 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=287 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=319 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=337 && yPixel<402) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=403 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=409 && yPixel<499) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=499 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=512 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=600 && yPixel<608) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=609 && yPixel<622) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=622 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=0 && xPixel<1 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=0 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=126 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=145 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=252 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=271 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=273 && yPixel<275) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=276 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=287 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=312 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=319 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=336 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=402 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=409 && yPixel<498) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=498 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=516 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=606 && yPixel<621) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=621 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=1 && xPixel<2 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=0 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=124 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=126 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=134 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=147 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=250 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=287 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=292 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=320 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=338 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=408 && yPixel<493) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=493 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=521 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=606 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=616 && yPixel<622) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=2 && xPixel<3 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=0 && yPixel<125) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=126 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=134 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=146 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=249 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=290 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=317 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=339 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=403 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=407 && yPixel<492) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=492 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=498 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=518 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=521 && yPixel<557) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=557 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=561 && yPixel<598) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=601 && yPixel<606) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=606 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=3 && xPixel<4 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=0 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=126 && yPixel<127) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=132 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=139 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=146 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=250 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=296 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=317 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=339 && yPixel<490) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=490 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=502 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=517 && yPixel<555) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=555 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=563 && yPixel<598) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=598 && yPixel<606) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=606 && yPixel<611) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=612 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=624 && yPixel<629) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=629 && yPixel<635) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=4 && xPixel<5 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=0 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=132 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=145 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=152 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=251 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=295 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=316 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=339 && yPixel<489) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=491 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=497 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=502 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=516 && yPixel<556) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=556 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=563 && yPixel<598) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=611 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=627 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=5 && xPixel<6 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=0 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=130 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=152 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=251 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=294 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=317 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=337 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=343 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=364 && yPixel<488) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=500 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=516 && yPixel<555) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=555 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=563 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=609 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=623 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=6 && xPixel<7 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=0 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=153 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=252 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=295 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=308 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=316 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=340 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=344 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=360 && yPixel<385) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=390 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=495 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=500 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=506 && yPixel<553) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=553 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=562 && yPixel<602) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=605 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=610 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=614 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=7 && xPixel<8 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=0 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=156 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=249 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=252 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=262 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=300 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=312 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=349 && yPixel<357) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=359 && yPixel<362) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=362 && yPixel<382) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=390 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=487 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=496 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=498 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=502 && yPixel<517) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=518 && yPixel<553) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=553 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=563 && yPixel<572) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=575 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=580 && yPixel<584) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=584 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=588 && yPixel<602) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=602 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=606 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=8 && xPixel<9 && yPixel>=615 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=0 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=155 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=159 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=251 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=253 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=261 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=300 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=312 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=361 && yPixel<380) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=380 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=383 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=390 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=487 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=494 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=499 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=516 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=521 && yPixel<552) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=552 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=567 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=600 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=605 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=9 && xPixel<10 && yPixel>=616 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=0 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=153 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=158 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=253 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=261 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=300 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=309 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=360 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=389 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=403 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=487 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=492 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=497 && yPixel<517) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=518 && yPixel<521) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=522 && yPixel<525) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=525 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=528 && yPixel<543) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=549 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=560 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=592 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=605 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=10 && xPixel<11 && yPixel>=616 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=0 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=159 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=254 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=257 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=260 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=298 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=302 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=311 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=352 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=359 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=385 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=388 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=403 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=441 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=496 && yPixel<525) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=525 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=532 && yPixel<539) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=539 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=553 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=558 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=569 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=575 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=585 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=592 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=604 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=615 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=11 && xPixel<12 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=0 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=151 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=201 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=204 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=255 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=303 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=311 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=356 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=377 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=381 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=385 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=403 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=440 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=442 && yPixel<482) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=484 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=495 && yPixel<525) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=525 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=551 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=574 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=584 && yPixel<591) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=592 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=604 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=614 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=12 && xPixel<13 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=0 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=205 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=252 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=303 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=311 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=351 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=356 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=361 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=377 && yPixel<380) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=381 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=384 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=403 && yPixel<419) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=420 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=441 && yPixel<483) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=496 && yPixel<520) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=524 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=545 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=570 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=593 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=604 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=618 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=13 && xPixel<14 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=0 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=200 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=206 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=251 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=303 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=310 && yPixel<353) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=353 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=356 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=376 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=383 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=398 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=402 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=411 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=415 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=431 && yPixel<484) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=484 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=494 && yPixel<517) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=519 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=544 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=563 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=592 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=605 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=14 && xPixel<15 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=0 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=196 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=206 && yPixel<248) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=249 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=297 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=304 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=355 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=375 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=383 && yPixel<394) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=394 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=401 && yPixel<410) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=415 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=431 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=495 && yPixel<517) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=517 && yPixel<529) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=530 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=541 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=15 && xPixel<16 && yPixel>=601 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=0 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=194 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=202 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=205 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=245 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=287 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=293 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=306 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=354 && yPixel<382) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=383 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=394 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=397 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=415 && yPixel<428) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=431 && yPixel<483) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=485 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=495 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=516 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=527 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=538 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=563 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=574 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=579 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=16 && xPixel<17 && yPixel>=600 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=0 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=194 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=202 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=205 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=245 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=285 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=290 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=304 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=341 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=347 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=352 && yPixel<378) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=380 && yPixel<391) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=392 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=396 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=410 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=415 && yPixel<427) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=427 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=433 && yPixel<483) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=484 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=487 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=492 && yPixel<515) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=515 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=532 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=563 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=575 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=588 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=599 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=633 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=17 && xPixel<18 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=0 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=194 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=202 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=205 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=244 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=285 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=304 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=348 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=352 && yPixel<361) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=365 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=380 && yPixel<390) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=392 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=397 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=402 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=406 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=415 && yPixel<425) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=432 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=445 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=453 && yPixel<484) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=484 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=486 && yPixel<488) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=492 && yPixel<509) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=509 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=526 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=563 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=573 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=588 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=599 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=18 && xPixel<19 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=0 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=153 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=191 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=202 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=204 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=244 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=285 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=310 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=341 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=351 && yPixel<361) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=361 && yPixel<367) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=367 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=379 && yPixel<388) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=388 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=393 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=414 && yPixel<422) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=422 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=428 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=432 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=444 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=454 && yPixel<488) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=491 && yPixel<507) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=507 && yPixel<520) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=520 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=561 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=574 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=592 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=19 && xPixel<20 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=0 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=101 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=153 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=191 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=202 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=204 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=242 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=284 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=312 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=333 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=342 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=357 && yPixel<362) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=362 && yPixel<365) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=367 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=378 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=388 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=390 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=414 && yPixel<422) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=424 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=428 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=432 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=445 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=451 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=454 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=491 && yPixel<505) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=505 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=518 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=576 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=629 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=20 && xPixel<21 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=0 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=76 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=93 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=101 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=151 && yPixel<189) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=189 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=192 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=204 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=241 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=284 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=309 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=313 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=342 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=347 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=349 && yPixel<353) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=353 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=358 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=389 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=416 && yPixel<421) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=421 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=431 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=444 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=454 && yPixel<486) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=491 && yPixel<503) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=503 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=518 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=574 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=628 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=21 && xPixel<22 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=0 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=102 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=147 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=153 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=192 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=201 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=239 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=284 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=303 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=313 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=317 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=344 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=356 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=386 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=400 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=404 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=417 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=420 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=427 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=434 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=446 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=449 && yPixel<451) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=455 && yPixel<458) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=459 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=487 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=492 && yPixel<499) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=499 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=513 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=576 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=22 && xPixel<23 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=0 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=90 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=93 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=99 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=152 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=190 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=201 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=239 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=285 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=302 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=304 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=319 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=349 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=357 && yPixel<388) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=388 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=394 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=395 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=399 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=405 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=417 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=420 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=431 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=437 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=447 && yPixel<449) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=449 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=462 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=487 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=493 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=512 && yPixel<542) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=546 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=578 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=632 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=23 && xPixel<24 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=0 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=80 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=98 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=146 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=152 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=190 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=195 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=200 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=238 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=285 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=300 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=305 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=313 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=322 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=347 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=355 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=387 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=392 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=396 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=405 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=415 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=419 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=437 && yPixel<448) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=451 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=462 && yPixel<486) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=486 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=491 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=496 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=498 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=502 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=506 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=541 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=547 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=578 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=24 && xPixel<25 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=0 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=100 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=147 && yPixel<189) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=190 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=199 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=235 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=284 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=300 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=305 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=319 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=354 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=387 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=390 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=397 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=399 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=402 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=413 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=420 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=437 && yPixel<448) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=459 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=464 && yPixel<484) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=484 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=490 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=500 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=502 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=505 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=510 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=538 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=549 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=567 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=578 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=588 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=25 && xPixel<26 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=0 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=96 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=152 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=198 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=234 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=284 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=299 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=305 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=319 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=352 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=391 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=406 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=413 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=423 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=438 && yPixel<447) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=447 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=452 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=459 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=465 && yPixel<483) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=483 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=492 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=496 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=502 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=536 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=549 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=565 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=26 && xPixel<27 && yPixel>=588 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=0 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=147 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=234 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=284 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=299 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=309 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=313 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=341 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=352 && yPixel<385) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=389 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=403 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=413 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=424 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=430 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=436 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=439 && yPixel<446) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=452 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=462 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=466 && yPixel<480) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=480 && yPixel<485) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=485 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=498 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=509 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=535 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=549 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=562 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=582 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=27 && xPixel<28 && yPixel>=589 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=0 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=147 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=152 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=195 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=234 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=284 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=300 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=313 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=344 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=351 && yPixel<385) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=386 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=402 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=409 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=414 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=431 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=436 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=439 && yPixel<446) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=446 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=450 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=453 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=464 && yPixel<484) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=484 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=492 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=499 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=509 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=534 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=542 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=548 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=558 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=565 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=590 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=28 && xPixel<29 && yPixel>=601 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=0 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=151 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=196 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=231 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=233 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=284 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=298 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=307 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=311 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=336 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=345 && yPixel<385) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=387 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=394 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=400 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=407 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=415 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=425 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=431 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=436 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=445 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=451 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=466 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=471 && yPixel<473) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=473 && yPixel<481) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=481 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=494 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=535 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=541 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=551 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=558 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=562 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=590 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=602 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=29 && xPixel<30 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=0 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=147 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=196 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=231 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=285 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=295 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=311 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=337 && yPixel<390) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=390 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=394 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=405 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=421 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=427 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=431 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=439 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=443 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=449 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=468 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=469 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=492 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=538 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=550 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=594 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=606 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=30 && xPixel<31 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=0 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=194 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=201 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=231 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=284 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=295 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=336 && yPixel<378) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=402 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=420 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=425 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=429 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=433 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=444 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=449 && yPixel<485) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=492 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=538 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=549 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=595 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=31 && xPixel<32 && yPixel>=616 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=0 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=193 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=198 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=231 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=292 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=336 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=378 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=383 && yPixel<390) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=402 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=412 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=418 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=422 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=432 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=447 && yPixel<485) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=487 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=492 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=533 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=539 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=550 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=597 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=32 && xPixel<33 && yPixel>=615 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=0 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=197 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=230 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=291 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=325 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=336 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=376 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=382 && yPixel<390) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=410 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=415 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=430 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=446 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=486 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=490 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=535 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=550 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=598 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=612 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=33 && xPixel<34 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=0 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=191 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=195 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=229 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=336 && yPixel<375) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=375 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=381 && yPixel<390) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=391 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=404 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=410 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=414 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=422 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=429 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=454 && yPixel<485) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=490 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=605 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=609 && yPixel<637) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=34 && xPixel<35 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=0 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=226 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=229 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=337 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=345 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=374 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=380 && yPixel<402) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=404 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=410 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=416 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=425 && yPixel<428) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=428 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=433 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=440 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=448 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=451 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=467 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=475 && yPixel<481) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=482 && yPixel<485) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=486 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=541 && yPixel<637) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=35 && xPixel<36 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=0 && yPixel<226) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=226 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=341 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=373 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=379 && yPixel<403) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=403 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=406 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=428 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=445 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=450 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=472 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=474 && yPixel<476) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=476 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=537 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=36 && xPixel<37 && yPixel>=541 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=0 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=105 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=227 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=335 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=342 && yPixel<372) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=373 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=378 && yPixel<404) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=407 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=422 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=425 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=445 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=448 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=471 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=535 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=541 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=574 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=37 && xPixel<38 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=0 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=224 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=282 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=342 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=373 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=377 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=415 && yPixel<421) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=424 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=430 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=434 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=445 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=465 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=468 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=470 && yPixel<472) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=472 && yPixel<475) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=475 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=536 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=539 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=549 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=559 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=569 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=38 && xPixel<39 && yPixel>=575 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=0 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=98 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=105 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=223 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=262 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=281 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=341 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=375 && yPixel<398) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=400 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=422 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=440 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=466 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=548 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=567 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=576 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=627 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=39 && xPixel<40 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=0 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=104 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=106 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=222 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=262 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=264 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=279 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=339 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=343 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=355 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=397 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=401 && yPixel<410) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=414 && yPixel<419) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=422 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=427 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=432 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=435 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=438 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=546 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=577 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=625 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=40 && xPixel<41 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=0 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=223 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=235 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=245 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=256 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=266 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=282 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=340 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=348 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=356 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=397 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=403 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=407 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=418 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=424 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=444 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=452 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=464 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=546 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=574 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=626 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=41 && xPixel<42 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=0 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=221 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=236 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=245 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=253 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=265 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=268 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=281 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=342 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=351 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=359 && yPixel<396) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=398 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=403 && yPixel<406) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=416 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=423 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=429 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=441 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=456 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=462 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=545 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=556 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=573 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=624 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=634 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=42 && xPixel<43 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=0 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=221 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=237 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=242 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=246 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=254 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=281 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=359 && yPixel<394) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=396 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=406 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=418 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=430 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=435 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=440 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=447 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=462 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=545 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=571 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=623 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=43 && xPixel<44 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=0 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=222 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=228 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=242 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=247 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=254 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=272 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=279 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=349 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=353 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=360 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=393 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=399 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=411 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=416 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=432 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=438 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=454 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=458 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=462 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=546 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=570 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=617 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=626 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=44 && xPixel<45 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=0 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=221 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=229 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=243 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=248 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=256 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=270 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=277 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=353 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=359 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=395 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=400 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=406 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=418 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=423 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=441 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=456 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=547 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=571 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=45 && xPixel<46 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=0 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=220 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=248 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=258 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=271 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=279 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=349 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=359 && yPixel<366) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=370 && yPixel<391) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=404 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=407 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=415 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=427 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=440 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=454 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=550 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=571 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=623 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=628 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=46 && xPixel<47 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=0 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=219 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=247 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=258 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=279 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=283 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=349 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=363 && yPixel<368) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=376 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=391 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=403 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=421 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=448 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=552 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=571 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=610 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=621 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=628 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=47 && xPixel<48 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=0 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=219 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=255 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=257 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=284 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=343 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=347 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=358 && yPixel<363) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=377 && yPixel<388) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=388 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=403 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=415 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=421 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=438 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=443 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=553 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=571 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=608 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=621 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=48 && xPixel<49 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=0 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=219 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=252 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=256 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=287 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=335 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=358 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=373 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=377 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=387 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=422 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=442 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=553 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=571 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=603 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=49 && xPixel<50 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=0 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=217 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=220 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=252 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=256 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=275 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=279 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=283 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=285 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=333 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=359 && yPixel<371) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=371 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=377 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=388 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=400 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=404 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=410 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=422 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=440 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=553 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=570 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=599 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=50 && xPixel<51 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=0 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=218 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=224 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=230 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=256 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=285 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=333 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=360 && yPixel<367) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=367 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=371 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=375 && yPixel<378) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=378 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=386 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=395 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=402 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=416 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=419 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=439 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=511 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=519 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=537 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=540 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=553 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=574 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=597 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=629 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=51 && xPixel<52 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=0 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=219 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=222 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=229 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=233 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=256 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=285 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=333 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=363 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=369 && yPixel<371) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=371 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=377 && yPixel<385) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=388 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=405 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=412 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=419 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=437 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=509 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=512 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=516 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=518 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=540 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=553 && yPixel<581) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=593 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=626 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=632 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=52 && xPixel<53 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=0 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=224 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=230 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=254 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=285 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=336 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=360 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=369 && yPixel<372) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=377 && yPixel<384) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=387 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=403 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=418 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=422 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=437 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=508 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=512 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=519 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=538 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=555 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=573 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=581 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=589 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=616 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=624 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=53 && xPixel<54 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=2 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=225 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=229 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=254 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=286 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=336 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=359 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=371 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=377 && yPixel<383) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=386 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=405 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=414 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=505 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=508 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=512 && yPixel<520) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=520 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=555 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=580 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=589 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=611 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=621 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=54 && xPixel<55 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=3 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=228 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=251 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=254 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=286 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=333 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=376 && yPixel<380) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=383 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=385 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=415 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=425 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=437 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=504 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=510 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=521 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=566 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=579 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=588 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=604 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=610 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=628 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=55 && xPixel<56 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=3 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=55 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=224 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=247 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=251 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=288 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=334 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=362 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=364 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=380 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=384 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=394 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=407 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=413 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=420 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=425 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=436 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=448 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=510 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=519 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=567 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=578 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=600 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=605 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=609 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=56 && xPixel<57 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=1 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=3 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=52 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=59 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=222 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=246 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=256 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=263 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=289 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=334 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=362 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=364 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=401 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=406 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=417 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=421 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=425 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=429 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=436 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=448 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=513 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=518 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=567 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=578 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=608 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=57 && xPixel<58 && yPixel>=622 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=4 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=49 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=60 && yPixel<181) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=182 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=223 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=243 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=263 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=288 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=334 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=390 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=400 && yPixel<413) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=413 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=419 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=434 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=452 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=512 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=569 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=577 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=58 && xPixel<59 && yPixel>=619 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=1 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=4 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=46 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=63 && yPixel<172) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=179 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=219 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=232 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=241 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=263 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=287 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=302 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=333 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=360 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=391 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=397 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=399 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=413 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=420 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=435 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=444 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=514 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=559 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=615 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=59 && xPixel<60 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=7 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=42 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=50 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=56 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=64 && yPixel<181) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=182 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=222 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=238 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=266 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=289 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=300 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=306 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=331 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=352 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=361 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=389 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=395 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=414 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=424 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=430 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=446 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=560 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=613 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=634 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=60 && xPixel<61 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=4 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=6 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=9 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=11 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=20 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=46 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=50 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=57 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=63 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=223 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=241 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=266 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=289 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=298 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=305 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=311 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=330 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=351 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=353 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=361 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=393 && yPixel<409) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=409 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=417 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=429 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=446 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=455 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=466 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=560 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=603 && yPixel<613) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=615 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=632 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=61 && xPixel<62 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=4 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=6 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=12 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=15 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=18 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=46 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=50 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=63 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=240 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=261 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=265 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=292 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=315 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=322 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=328 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=351 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=353 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=361 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=389 && yPixel<409) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=409 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=452 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=455 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=561 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=573 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=601 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=616 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=62 && xPixel<63 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=9 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=15 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=18 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=46 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=51 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=62 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=259 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=264 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=289 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=321 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=352 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=361 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=389 && yPixel<408) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=411 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=416 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=449 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=451 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=456 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=573 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=584 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=599 && yPixel<613) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=615 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=63 && xPixel<64 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=9 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=12 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=17 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=39 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=47 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=51 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=62 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=264 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=290 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=320 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=361 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=389 && yPixel<408) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=412 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=450 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=457 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=564 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=571 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=600 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=609 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=64 && xPixel<65 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=8 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=13 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=16 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=40 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=44 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=46 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=49 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=61 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=259 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=266 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=287 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=289 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=318 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=361 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=385 && yPixel<388) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=389 && yPixel<403) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=409 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=414 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=459 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=560 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=571 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=583 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=604 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=65 && xPixel<66 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=7 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=9 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=12 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=15 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=17 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=43 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=46 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=61 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=263 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=291 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=318 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=352 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=360 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=389 && yPixel<402) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=404 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=409 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=414 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=464 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=561 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=571 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=579 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=584 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=596 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=630 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=66 && xPixel<67 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=5 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=7 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=17 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=39 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=43 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=61 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=231 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=293 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=318 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=352 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=358 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=387 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=394 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=397 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=409 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=415 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=442 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=447 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=450 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=468 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=562 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=578 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=584 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=621 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=628 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=67 && xPixel<68 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=13 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=18 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=39 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=61 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=233 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=293 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=318 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=344 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=352 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=358 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=388 && yPixel<395) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=395 && yPixel<398) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=402 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=413 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=418 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=430 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=440 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=443 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=449 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=466 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=494 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=562 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=573 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=579 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=584 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=591 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=618 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=627 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=68 && xPixel<69 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=8 && yPixel<16) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=19 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=40 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=61 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=288 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=293 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=314 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=317 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=344 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=352 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=355 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=359 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=396 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=412 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=420 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=424 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=428 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=452 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=468 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=499 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=574 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=584 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=606 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=613 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=69 && xPixel<70 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=13 && yPixel<16) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=19 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=38 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=42 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=61 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=287 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=293 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=313 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=316 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=344 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=352 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=358 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=405 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=423 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=447 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=452 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=468 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=495 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=500 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=576 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=583 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=605 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=70 && xPixel<71 && yPixel>=612 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=18 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=36 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=41 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=61 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=287 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=294 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=315 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=335 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=344 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=354 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=358 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=410 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=447 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=451 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=454 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=467 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=495 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=500 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=576 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=595 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=608 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=626 && yPixel<635) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=71 && xPixel<72 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=2 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=16 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=36 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=42 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=61 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=286 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=302 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=306 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=314 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=331 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=333 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=339 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=344 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=419 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=450 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=454 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=466 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=496 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=500 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=563 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=575 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=593 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=600 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=72 && xPixel<73 && yPixel>=625 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=1 && yPixel<6) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=6 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=9 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=12 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=34 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=43 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=58 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=60 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=283 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=312 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=318 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=344 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=424 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=449 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=454 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=463 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=467 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=497 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=500 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=562 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=575 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=600 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=73 && xPixel<74 && yPixel>=623 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=7 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=11 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=35 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=41 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=43 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=61 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=281 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=315 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=321 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=341 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=373 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=432 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=453 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=463 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=499 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=504 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=516 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=575 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=74 && xPixel<75 && yPixel>=623 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=2 && yPixel<7) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=7 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=12 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=34 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=41 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=45 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=62 && yPixel<275) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=275 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=306 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=321 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=380 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=437 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=441 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=452 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=461 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=501 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=505 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=513 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=515 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=567 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=575 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=75 && xPixel<76 && yPixel>=623 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=3 && yPixel<7) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=7 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=15 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=35 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=44 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=46 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=61 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=274 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=302 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=315 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=321 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=374 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=381 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=434 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=438 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=443 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=458 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=502 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=505 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=513 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=562 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=574 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=600 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=607 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=76 && xPixel<77 && yPixel>=623 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=4 && yPixel<8) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=8 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=16 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=34 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=45 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=60 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=269 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=272 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=301 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=313 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=322 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=335 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=359 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=374 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=381 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=416 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=419 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=437 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=445 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=560 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=570 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=598 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=609 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=77 && xPixel<78 && yPixel>=618 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=4 && yPixel<10) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=10 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=18 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=29 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=34 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=43 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=47 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=56 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=262 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=297 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=311 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=322 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=332 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=337 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=362 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=374 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=381 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=405 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=413 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=426 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=440 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=445 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=513 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=559 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=567 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=581 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=589 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=596 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=78 && xPixel<79 && yPixel>=621 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=5 && yPixel<9) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=9 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=19 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=33 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=42 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=55 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=261 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=297 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=308 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=322 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=328 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=337 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=346 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=356 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=362 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=369 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=374 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=381 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=405 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=411 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=445 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=569 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=579 && yPixel<594) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=79 && xPixel<80 && yPixel>=594 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=6 && yPixel<8) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=8 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=19 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=33 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=54 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=56 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=261 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=297 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=305 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=322 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=333 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=343 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=347 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=356 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=361 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=371 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=380 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=404 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=410 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=451 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=525 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=560 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=577 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=596 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=80 && xPixel<81 && yPixel>=615 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=24 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=35 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=56 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=261 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=296 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=312 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=323 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=332 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=347 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=360 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=367 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=376 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=380 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=409 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=434 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=443 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=451 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=454 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=516 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=528 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=560 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=573 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=586 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=81 && xPixel<82 && yPixel>=616 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=2 && yPixel<21) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=22 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=26 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=29 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=36 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=57 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=254 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=260 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=297 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=305 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=322 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=331 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=360 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=363 && yPixel<366) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=366 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=379 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=403 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=434 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=459 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=510 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=539 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=560 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=569 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=576 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=582 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=586 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=606 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=609 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=82 && xPixel<83 && yPixel>=616 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=22 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=30 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=33 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=39 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=58 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=87 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=252 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=255 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=261 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=299 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=306 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=315 && yPixel<325) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=325 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=337 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=356 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=362 && yPixel<366) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=376 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=378 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=400 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=433 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=462 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=508 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=513 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=524 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=541 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=551 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=561 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=568 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=573 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=586 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=83 && xPixel<84 && yPixel>=606 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=12 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=23 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=32 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=39 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=41 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=58 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=66 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=67 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=79 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=90 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=252 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=262 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=303 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=307 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=311 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=326 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=333 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=338 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=351 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=355 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=370 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=377 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=399 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=449 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=453 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=459 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=466 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=507 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=511 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=523 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=537 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=541 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=546 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=561 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=566 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=589 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=616 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=84 && xPixel<85 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=12 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=23 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=27 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=34 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=42 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=59 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=62 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=71 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=77 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=91 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=245 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=252 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=264 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=304 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=312 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=326 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=331 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=337 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=351 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=370 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=398 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=407 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=419 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=427 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=449 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=455 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=458 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=466 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=493 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=506 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=508 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=517 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=522 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=533 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=539 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=546 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=564 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=578 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=588 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=623 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=629 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=85 && xPixel<86 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=3 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=6 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=8 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=10 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=14 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=24 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=27 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=32 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=41 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=62 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=73 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=75 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=91 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=244 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=252 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=262 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=309 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=313 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=336 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=351 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=369 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=378 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=382 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=398 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=402 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=407 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=417 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=431 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=448 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=465 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=488 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=496 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=507 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=521 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=531 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=551 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=576 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=581 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=587 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=625 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=86 && xPixel<87 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=1 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=3 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=6 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=10 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=14 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=28 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=33 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=41 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=92 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=242 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=255 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=263 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=289 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=315 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=336 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=351 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=358 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=368 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=376 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=378 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=383 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=407 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=413 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=416 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=425 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=433 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=443 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=465 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=491 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=497 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=503 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=507 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=519 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=533 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=551 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=567 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=577 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=588 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=604 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=616 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=87 && xPixel<88 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=10 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=14 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=24 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=29 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=35 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=43 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=48 && yPixel<52) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=52 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=93 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=241 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=260 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=287 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=290 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=318 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=328 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=336 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=357 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=364 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=368 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=383 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=408 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=433 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=438 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=463 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=499 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=508 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=519 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=537 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=539 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=561 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=571 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=578 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=590 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=600 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=88 && xPixel<89 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=10 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=16 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=29 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=48 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=54 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=94 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=240 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=286 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=291 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=313 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=318 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=335 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=344 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=349 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=357 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=364 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=369 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=372 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=378 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=383 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=409 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=429 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=436 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=454 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=463 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=491 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=498 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=501 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=509 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=514 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=519 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=545 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=570 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=582 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=589 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=595 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=632 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=89 && xPixel<90 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=13 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=21 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=29 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=48 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=53 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=72 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=94 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=238 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=290 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=309 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=319 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=337 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=342 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=362 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=367 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=381 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=394 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=412 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=422 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=433 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=436 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=446 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=459 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=465 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=495 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=499 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=503 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=513 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=521 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=544 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=549 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=556 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=571 && yPixel<581) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=582 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=590 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=610 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=620 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=90 && xPixel<91 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=13 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=16 && yPixel<21) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=22 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=49 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=54 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=66 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=73 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=94 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=236 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=285 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=290 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=309 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=318 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=341 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=363 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=377 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=382 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=417 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=423 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=444 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=457 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=466 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=496 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=502 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=509 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=512 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=518 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=522 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=548 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=557 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=579 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=589 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=625 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=91 && xPixel<92 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=13 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=16 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=19 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=23 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=61 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=73 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=80 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=94 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=235 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=284 && yPixel<287) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=289 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=301 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=305 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=310 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=318 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=339 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=363 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=383 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=423 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=429 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=439 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=456 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=468 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=492 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=500 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=502 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=523 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=537 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=539 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=543 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=549 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=554 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=559 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=588 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=600 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=92 && xPixel<93 && yPixel>=622 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=14 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=27 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=30 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=61 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=69 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=80 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=95 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=239 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=288 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=306 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=310 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=320 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=335 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=363 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=371 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=383 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=417 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=423 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=428 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=435 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=437 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=455 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=462 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=491 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=503 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=516 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=524 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=534 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=545 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=558 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=583 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=588 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=608 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=623 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=93 && xPixel<94 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=15 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=32 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=52 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=54 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=62 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=69 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=78 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=79 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=96 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=241 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=243 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=302 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=310 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=320 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=327 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=94 && xPixel<95 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=94 && xPixel<95 && yPixel>=344 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=354 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=94 && xPixel<95 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=360 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=371 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=383 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=417 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=431 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=460 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=487 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=493 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=503 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=513 && yPixel<530) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=533 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=584 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=588 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=621 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=94 && xPixel<95 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=0 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=16 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=20 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=25 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=31 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=50 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=55 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=69 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=95 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=251 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=306 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=328 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=338 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b11000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=95 && xPixel<96 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=377 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=382 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=401 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=417 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=426 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=457 && yPixel<485) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=485 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=493 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=503 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=507 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=533 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=542 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=551 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=579 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=584 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=587 && yPixel<591) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=591 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=629 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=95 && xPixel<96 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=0 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=30 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=48 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=56 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=73 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=76 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=92 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=95 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=106 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=109 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=110 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=113 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=251 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=253 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=317 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=336 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b11000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b11000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=96 && xPixel<97 && yPixel>=351 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=360 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=366 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=381 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=401 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=423 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=455 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=458 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=483 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=492 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=534 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=539 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=553 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=579 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=588 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=599 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=615 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=626 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=96 && xPixel<97 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=0 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=36 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=49 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=57 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=62 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=65 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=74 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=76 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=87 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=98 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=105 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=115 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=117 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=118 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=119 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=120 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=254 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=296 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=320 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=334 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=97 && xPixel<98 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b11000000,8'b11111111};
	if(xPixel>=97 && xPixel<98 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=97 && xPixel<98 && yPixel>=342 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=97 && xPixel<98 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=351 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=359 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=381 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=385 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=388 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=416 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=433 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=452 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=456 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=483 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=490 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=562 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=579 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=589 && yPixel<591) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=595 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=612 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=627 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=97 && xPixel<98 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=0 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=37 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=58 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=63 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=66 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=67 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=76 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=102 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=104 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=122 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=255 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=295 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=305 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=313 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=323 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=98 && xPixel<99 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b11000000,8'b11111111};
	if(xPixel>=98 && xPixel<99 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=98 && xPixel<99 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=98 && xPixel<99 && yPixel>=340 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=350 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=391 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=412 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=420 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=434 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=450 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=457 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=487 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=518 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=521 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=536 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=567 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=578 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=590 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=623 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=98 && xPixel<99 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=7 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=23 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=38 && yPixel<50) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=50 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=57 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=65 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=71 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=75 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=123 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=126 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=253 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=256 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=277 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=295 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=303 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=323 && yPixel<327) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=327 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=340 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=365 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=377 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=383 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=390 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=410 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=427 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=431 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=433 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=438 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=443 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=451 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=456 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=516 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=521 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=537 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=578 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=589 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=617 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=629 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=99 && xPixel<100 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=2 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=4 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=7 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=13 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=22 && yPixel<26) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=26 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=38 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=49 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=72 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=124 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=128 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=137 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=138 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=255 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=292 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=302 && yPixel<325) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=329 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=340 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=347 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=357 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=368 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=375 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=380 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=383 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=387 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=390 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=410 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=426 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=439 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=443 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=456 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=519 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=535 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=540 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=568 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=572 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=585 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=610 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=628 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=633 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=100 && xPixel<101 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=4 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=7 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=13 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=20 && yPixel<28) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=28 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=39 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=49 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=52 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=61 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=73 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=115 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=125 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=133 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=137 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=138 && yPixel<143) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=143 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=147 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=153 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=255 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=279 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=288 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=302 && yPixel<327) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=346 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=356 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=368 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=390 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=399 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=404 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=407 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=420 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=431 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=435 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=441 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=445 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=457 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=515 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=517 && yPixel<530) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=530 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=541 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=572 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=582 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=585 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=608 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=615 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=623 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=633 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=101 && xPixel<102 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=1 && yPixel<2) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=2 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=13 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=20 && yPixel<48) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=48 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=53 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=63 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=72 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=87 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=130 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=140 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=155 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=255 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=277 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=300 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=333 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=342 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=348 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=355 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=365 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=375 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=378 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=381 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=390 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=403 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=407 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=417 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=426 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=433 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=442 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=460 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=510 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=523 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=527 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=542 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=569 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=575 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=585 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=606 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=618 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=623 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=632 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=102 && xPixel<103 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=1 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=7 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=15 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=22 && yPixel<38) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=44 && yPixel<46) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=49 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=56 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=63 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=84 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=86 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=88 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=122 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=141 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=156 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=254 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=272 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=280 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=284 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=299 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=340 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=352 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=362 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=375 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=378 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=383 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=384 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=387 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=393 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=402 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=406 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=411 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=416 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=420 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=430 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=437 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=459 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=505 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=511 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=526 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=531 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=536 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=541 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=551 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=555 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=574 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=585 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=603 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=609 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=617 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=103 && xPixel<104 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=1 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=10 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=13 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=24 && yPixel<35) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=41 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=43 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=48 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=58 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=63 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=84 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=87 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=157 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=205 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=254 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=271 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=273 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=282 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=290 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=300 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=329 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=337 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=340 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=359 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=373 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=379 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=104 && xPixel<105 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=387 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=392 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=398 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=403 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=419 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=459 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=501 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=512 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=518 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=526 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=546 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=553 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=562 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=569 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=584 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=602 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=614 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=104 && xPixel<105 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=27 && yPixel<37) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=37 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=40 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=43 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=46 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=61 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=64 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=78 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=155 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=162 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=206 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=254 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=271 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=273 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=280 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=324 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=331 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=333 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=340 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=355 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=372 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=376 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=379 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=105 && xPixel<106 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=105 && xPixel<106 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=392 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=403 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=411 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=418 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=439 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=459 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=499 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=519 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=544 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=552 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=561 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=581 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=594 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=608 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=612 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=105 && xPixel<106 && yPixel>=625 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=8 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=31 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=34 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=39 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=54 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=62 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=64 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=144 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=150 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=156 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=160 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=163 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=206 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=256 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=273 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=283 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=322 && yPixel<325) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=325 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=344 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=349 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=353 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=371 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=376 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=106 && xPixel<107 && yPixel>=380 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=383 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=106 && xPixel<107 && yPixel>=384 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=106 && xPixel<107 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=106 && xPixel<107 && yPixel>=390 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=393 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=403 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=411 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=418 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=451 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=460 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=472 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=496 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=521 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=530 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=544 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=579 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=587 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=590 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=612 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=624 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=106 && xPixel<107 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=0 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=32 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=39 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=58 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=65 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=98 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=105 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=146 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=155 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=158 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=162 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=206 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=255 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=257 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=267 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=273 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=279 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=285 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=327 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=331 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=335 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=344 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=353 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=370 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=373 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=378 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=107 && xPixel<108 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=107 && xPixel<108 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=107 && xPixel<108 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=107 && xPixel<108 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=388 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=107 && xPixel<108 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=107 && xPixel<108 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=403 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=411 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=414 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=449 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=460 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=470 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=474 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=497 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=519 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=546 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=586 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=594 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=601 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=607 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=624 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=107 && xPixel<108 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=2 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=42 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=60 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=65 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=75 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=79 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=82 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=84 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=89 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=98 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=107 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=146 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=152 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=159 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=202 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=205 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=257 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=267 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=269 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=272 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=280 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=283 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=302 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=321 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=330 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=341 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=364 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=369 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=108 && xPixel<109 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=108 && xPixel<109 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=108 && xPixel<109 && yPixel>=376 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=108 && xPixel<109 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=401 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=413 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=440 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=447 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=461 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=473 && yPixel<479) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=481 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=497 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=519 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=547 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=570 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=575 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=580 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=592 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=613 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=619 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=108 && xPixel<109 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=3 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=42 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=60 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=64 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=73 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=80 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=83 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=87 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=90 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=102 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=107 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=152 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=158 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=199 && yPixel<205) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=206 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=257 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=269 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=272 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=288 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=294 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=303 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=321 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=358 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=370 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=373 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=109 && xPixel<110 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=401 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=408 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=412 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=422 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=434 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=451 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=460 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=467 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=473 && yPixel<477) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=478 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=496 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=519 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=540 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=546 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=574 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=577 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=607 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=614 && yPixel<637) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=109 && xPixel<110 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=6 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=45 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=64 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=74 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=84 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=91 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=95 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=99 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=159 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=198 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=206 && yPixel<211) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=212 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=256 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=266 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=272 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=298 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=320 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=357 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=110 && xPixel<111 && yPixel>=371 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=110 && xPixel<111 && yPixel>=390 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=393 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=400 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=409 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=413 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=421 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=445 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=453 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=461 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=467 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=471 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=474 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=496 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=518 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=544 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=568 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=575 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=596 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=604 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=613 && yPixel<622) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=624 && yPixel<635) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=110 && xPixel<111 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=6 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=46 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=62 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=75 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=82 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=93 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=99 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=159 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=199 && yPixel<208) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=211 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=216 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=256 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=269 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=274 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=319 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=323 && yPixel<325) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=325 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=335 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=359 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=367 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=369 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=111 && xPixel<112 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=111 && xPixel<112 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=393 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=400 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=404 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=413 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=420 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=445 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=454 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=461 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=472 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=500 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=502 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=517 && yPixel<520) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=520 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=527 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=543 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=559 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=574 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=591 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=596 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=602 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=619 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=624 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=628 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=111 && xPixel<112 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=5 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=9 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=14 && yPixel<18) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=18 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=46 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=58 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=76 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=78 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=87 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=98 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=120 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=125 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=160 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=198 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=207 && yPixel<212) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=216 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=222 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=229 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=255 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=265 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=268 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=274 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=299 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=304 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=312 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=318 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=323 && yPixel<325) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=330 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=338 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=112 && xPixel<113 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=358 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=112 && xPixel<113 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=112 && xPixel<113 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=112 && xPixel<113 && yPixel>=369 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=112 && xPixel<113 && yPixel>=373 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=112 && xPixel<113 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=393 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=405 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=412 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=420 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=458 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=470 && yPixel<479) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=481 && yPixel<484) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=490 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=502 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=518 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=528 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=540 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=550 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=572 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=586 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=597 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=613 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=624 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=628 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=112 && xPixel<113 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=6 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=9 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=14 && yPixel<21) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=21 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=47 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=57 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=62 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=68 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=71 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=82 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=87 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=91 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=121 && yPixel<131) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=131 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=164 && yPixel<179) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=179 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=188 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=195 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=206 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=216 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=223 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=243 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=246 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=255 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=265 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=272 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=299 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=304 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=315 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=321 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=328 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=340 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=348 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=352 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=359 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=113 && xPixel<114 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=372 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=113 && xPixel<114 && yPixel>=388 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=394 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=400 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=404 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=421 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=466 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=469 && yPixel<477) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=477 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=489 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=502 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=509 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=512 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=518 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=522 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=527 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=539 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=569 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=581 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=595 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=600 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=626 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=113 && xPixel<114 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=7 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=10 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=19 && yPixel<22) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=22 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=47 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=57 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=62 && yPixel<67) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=67 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=71 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=81 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=87 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=94 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=123 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=125 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=164 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=170 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=179 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=186 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=188 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=195 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=206 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=220 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=246 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=254 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=290 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=297 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=304 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=307 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=314 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=323 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=329 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=340 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=344 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=353 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=114 && xPixel<115 && yPixel>=359 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=114 && xPixel<115 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=114 && xPixel<115 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=114 && xPixel<115 && yPixel>=368 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=114 && xPixel<115 && yPixel>=372 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=114 && xPixel<115 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=395 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=403 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=416 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=420 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=467 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=474 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=489 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=498 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=503 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=514 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=524 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=538 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=544 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=566 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=579 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=584 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=593 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=598 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=615 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=623 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=114 && xPixel<115 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=10 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=27 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=49 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=55 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=62 && yPixel<67) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=67 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=71 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=75 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=95 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=108 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=140 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=174 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=180 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=191 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=198 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=206 && yPixel<211) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=211 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=219 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=254 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=294 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=299 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=305 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=323 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=328 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=340 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=344 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=348 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=354 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=115 && xPixel<116 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=115 && xPixel<116 && yPixel>=373 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=115 && xPixel<116 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=115 && xPixel<116 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=390 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=402 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=409 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=462 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=466 && yPixel<472) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=472 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=489 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=499 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=510 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=515 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=520 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=527 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=536 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=544 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=562 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=569 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=572 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=580 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=597 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=612 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=622 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=115 && xPixel<116 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=11 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=27 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=49 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=56 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=62 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=68 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=72 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=87 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=88 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=96 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=105 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=113 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=139 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=144 && yPixel<156) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=156 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=180 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=190 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=195 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=198 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=204 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=217 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=254 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=280 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=292 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=300 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=305 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=314 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=321 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=327 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=332 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=340 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=347 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=356 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=362 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=365 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=367 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=116 && xPixel<117 && yPixel>=376 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11111111};
	if(xPixel>=116 && xPixel<117 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=382 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=388 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=402 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=407 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=461 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=465 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=471 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=495 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=503 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=508 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=513 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=520 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=528 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=532 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=558 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=563 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=570 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=597 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=608 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=617 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=622 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=116 && xPixel<117 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=8 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=12 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=50 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=56 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=62 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=66 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=72 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=87 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=106 && yPixel<127) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=127 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=138 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=144 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=160 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=179 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=192 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=199 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=210 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=216 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=256 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=273 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=277 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=283 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=301 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=117 && xPixel<118 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=320 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=327 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=333 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=340 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=357 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11111111};
	if(xPixel>=117 && xPixel<118 && yPixel>=373 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=383 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=386 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=400 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=405 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=459 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=464 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=468 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=491 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=499 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=512 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=515 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=518 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=523 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=527 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=569 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=594 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=605 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=629 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=117 && xPixel<118 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=7 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=12 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=50 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=56 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=62 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=66 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=73 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=83 && yPixel<88) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=88 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=106 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=141 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=145 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=162 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=178 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=191 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=193 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=197 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=215 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=254 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=257 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=273 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=283 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=301 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=311 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=118 && xPixel<119 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b11000000,8'b11111111};
	if(xPixel>=118 && xPixel<119 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=118 && xPixel<119 && yPixel>=317 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=333 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=340 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=342 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=358 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=366 && yPixel<369) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=369 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=384 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=395 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=399 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=404 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=457 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=464 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=493 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=497 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=512 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=516 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=519 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=559 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=585 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=606 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=618 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=627 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=118 && xPixel<119 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=6 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=13 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=48 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=56 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=73 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=80 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=83 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=90 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=107 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=157 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=161 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=176 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=192 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=197 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=200 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=216 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=235 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=259 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=273 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=282 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=306 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11111111};
	if(xPixel>=119 && xPixel<120 && yPixel>=316 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=329 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=335 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=341 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=368 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=382 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=393 && yPixel<397) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=398 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=455 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=463 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=488 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=495 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=507 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=516 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=546 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=550 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=563 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=581 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=597 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=605 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=612 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=618 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=119 && xPixel<120 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=2 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=4 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=9 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=13 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=28 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=49 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=57 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=73 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=78 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=83 && yPixel<88) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=88 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=92 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=108 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=125 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=132 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=150 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=158 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=175 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=201 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=218 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=260 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=273 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=281 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=305 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=329 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=340 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=342 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=378 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=391 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=397 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=454 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=460 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=493 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=499 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=502 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=516 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=551 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=558 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=565 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=581 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=590 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=597 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=610 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=615 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=621 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=120 && xPixel<121 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=1 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=2 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=25 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=28 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=49 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=59 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=73 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=75 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=82 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=92 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=116 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=119 && yPixel<124) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=124 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=132 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=139 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=147 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=158 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=175 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=203 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=218 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=221 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=227 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=237 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=260 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=272 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=279 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=298 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=305 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=326 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=333 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=345 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=396 && yPixel<416) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=417 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=452 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=481 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=486 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=495 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=500 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=510 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=516 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=519 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=548 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=553 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=577 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=595 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=611 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=624 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=121 && xPixel<122 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=28 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=51 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=57 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=61 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=74 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=77 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=81 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=90 && yPixel<92) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=93 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=137 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=141 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=148 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=161 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=169 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=176 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=216 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=231 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=236 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=272 && yPixel<275) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=278 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=284 && yPixel<287) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=287 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=297 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=305 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=339 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=345 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=380 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=391 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=394 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=419 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=435 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=450 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=460 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=477 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=479 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=484 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=497 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=500 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=503 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=511 && yPixel<520) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=520 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=568 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=582 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=611 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=625 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=122 && xPixel<123 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=0 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=28 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=31 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=51 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=59 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=65 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=73 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=76 && yPixel<78) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=78 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=83 && yPixel<88) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=88 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=90 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=95 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=121 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=157 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=170 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=174 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=217 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=229 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=232 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=263 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=288 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=298 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=305 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=313 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=332 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=335 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=367 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=388 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=393 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=414 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=429 && yPixel<436) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=439 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=448 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=492 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=498 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=514 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=522 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=551 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=556 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=560 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=576 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=580 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=608 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=615 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=625 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=123 && xPixel<124 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=1 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=4 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=15 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=28 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=33 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=51 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=68 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=73 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=82 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=89 && yPixel<92) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=94 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=99 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=105 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=108 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=109 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=118 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=125 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=149 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=157 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=173 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=223 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=229 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=232 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=263 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=276 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=314 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=318 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=328 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=334 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=359 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=370 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=386 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=392 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=414 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=431 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=439 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=446 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=490 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=500 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=506 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=509 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=511 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=514 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=522 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=542 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=568 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=594 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=610 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=124 && xPixel<125 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=1 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=2 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=3 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=5 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=29 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=34 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=54 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=67 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=73 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=77 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=80 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=84 && yPixel<86) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=87 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=90 && yPixel<92) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=95 && yPixel<100) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=100 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=104 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=108 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=116 && yPixel<128) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=128 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=139 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=157 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=172 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=223 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=231 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=276 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=305 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=320 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=334 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=358 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=372 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=386 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=391 && yPixel<412) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=412 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=444 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=485 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=489 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=496 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=506 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=510 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=516 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=521 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=537 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=567 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=600 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=608 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=613 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=623 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=125 && xPixel<126 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=4 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=6 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=31 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=36 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=54 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=66 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=73 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=77 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=80 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=87 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=99 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=104 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=107 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=113 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=118 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=119 && yPixel<128) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=128 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=137 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=151 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=157 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=172 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=222 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=230 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=276 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=291 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=300 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=306 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=324 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=332 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=354 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=378 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=385 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=388 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=403 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=415 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=442 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=458 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=469 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=475 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=484 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=490 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=509 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=516 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=519 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=536 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=545 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=568 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=589 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=596 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=601 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=609 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=614 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=623 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=126 && xPixel<127 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=5 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=7 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=53 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=66 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=70 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=73 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=77 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=85 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=93 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=96 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=101 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=104 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=107 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=111 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=122 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=125 && yPixel<127) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=127 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=137 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=145 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=157 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=165 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=172 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=179 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=185 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=190 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=217 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=229 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=276 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=282 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=289 && yPixel<300) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=302 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=311 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=322 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b11000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=337 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=352 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=384 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=387 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=402 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=410 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=440 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=456 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=474 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=482 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=504 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=519 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=533 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=536 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=545 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=570 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=594 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=605 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=611 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=619 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=624 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=127 && xPixel<128 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=7 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=10 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=53 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=57 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=65 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=69 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=73 && yPixel<76) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=76 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=91 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=98 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=100 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=104 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=107 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=112 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=118 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=132 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=139 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=169 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=171 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=178 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=182 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=190 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=215 && yPixel<226) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=229 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=263 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=272 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=287 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=305 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=313 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=349 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=386 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=410 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=438 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=453 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=476 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=481 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=505 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=516 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=519 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=530 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=532 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=545 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=571 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=584 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=590 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=594 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=605 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=609 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b11000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=627 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=633 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=128 && xPixel<129 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=7 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=9 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=12 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=47 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=57 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=61 && yPixel<63) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=63 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=73 && yPixel<76) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=76 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=79 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=86 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=92 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=97 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=105 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=107 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=112 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=116 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=121 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=141 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=173 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=177 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=183 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=197 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=214 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=227 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=261 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=287 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=313 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=347 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=380 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=385 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=405 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=408 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=431 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=436 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=448 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=474 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=484 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=489 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=508 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=517 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=533 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=545 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=572 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=580 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=604 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=609 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=623 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=630 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=129 && xPixel<130 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=6 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=12 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=39 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=42 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=48 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=60 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=82 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=86 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=99 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=102 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=105 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=111 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=115 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=119 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=120 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=140 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=153 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=172 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=177 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=183 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=199 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=213 && yPixel<222) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=225 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=261 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=281 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=287 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=312 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=319 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=329 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=346 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=379 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=384 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=395 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=409 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=433 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=436 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=472 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=475 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=481 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=508 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=516 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=533 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=545 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=552 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=562 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=570 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=576 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=591 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=595 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=609 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=622 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=628 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=130 && xPixel<131 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=5 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=11 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=42 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=61 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=69 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=81 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=85 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=104 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=110 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=113 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=137 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=151 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=155 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=161 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=186 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=193 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=200 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=216 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=220 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=261 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=266 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=281 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=287 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=311 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=320 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=333 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=378 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=382 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=392 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=402 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=409 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=427 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=433 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=463 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=470 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=472 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=476 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=484 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=515 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=517 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=531 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=534 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=548 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=555 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=575 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=583 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=589 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=616 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=620 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=131 && xPixel<132 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=8 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=11 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=41 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=49 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=62 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=64 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=74 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=89 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=110 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=112 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=122 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=126 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=136 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=145 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=165 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=177 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=186 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=200 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=214 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=220 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=263 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=272 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=276 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=281 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=288 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=310 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=323 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=335 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=378 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=381 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=391 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=400 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=406 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=409 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=425 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=431 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=461 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=470 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=473 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=513 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=519 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=539 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=577 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=590 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=624 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=132 && xPixel<133 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=11 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=44 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=52 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=56 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=63 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=74 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=81 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=87 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=105 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=110 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=115 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=118 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=126 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=135 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=146 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=162 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=169 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=185 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=188 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=200 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=214 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=220 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=258 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=263 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=266 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=270 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=274 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=279 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=288 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=310 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=322 && yPixel<325) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=325 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=335 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=375 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=381 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=391 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=399 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=413 && yPixel<417) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=417 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=423 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=428 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=466 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=471 && yPixel<478) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=478 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=481 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=514 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=519 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=561 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=577 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=585 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=592 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=624 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=632 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=133 && xPixel<134 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=14 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=43 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=52 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=72 && yPixel<78) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=81 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=89 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=112 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=116 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=119 && yPixel<123) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=123 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=126 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=131 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=135 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=144 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=160 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=186 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=202 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=219 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=242 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=252 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=256 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=265 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=269 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=273 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=282 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=291 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=310 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=324 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=335 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=351 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=364 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=382 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=391 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=396 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=405 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=418 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=424 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=469 && yPixel<476) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=476 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=487 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=491 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=507 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=514 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=520 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=530 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=574 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=586 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=595 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=619 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=627 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=134 && xPixel<135 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=15 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=43 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=45 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=47 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=50 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=72 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=75 && yPixel<78) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=81 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=95 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=112 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=114 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=116 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=118 && yPixel<124) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=124 && yPixel<127) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=127 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=131 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=140 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=160 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=170 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=182 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=201 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=219 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=241 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=245 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=251 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=255 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=261 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=270 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=292 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=309 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=323 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=338 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=346 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=350 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=364 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=373 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=379 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=384 && yPixel<391) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=391 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=396 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=405 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=416 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=422 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=463 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=466 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=468 && yPixel<475) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=476 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=480 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=490 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=504 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=518 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=525 && yPixel<539) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=539 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=578 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=594 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=598 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=605 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=626 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=135 && xPixel<136 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=12 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=16 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=43 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=51 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=77 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=82 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=99 && yPixel<102) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=102 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=112 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=119 && yPixel<123) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=123 && yPixel<128) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=130 && yPixel<132) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=133 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=139 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=163 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=166 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=177 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=183 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=195 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=205 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=220 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=239 && yPixel<248) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=249 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=254 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=260 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=265 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=268 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=274 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=292 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=310 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=322 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=336 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=343 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=353 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=360 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=371 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=377 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=393 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=400 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=406 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=417 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=466 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=474 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=481 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=488 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=494 && yPixel<502) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=502 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=525 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=532 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=537 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=540 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=576 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=580 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=594 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=611 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=619 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=136 && xPixel<137 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=0 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=16 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=45 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=54 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=69 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=76 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=79 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=85 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=89 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=93 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=99 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=106 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=112 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=115 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=118 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=122 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=126 && yPixel<131) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=131 && yPixel<135) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=137 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=142 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=160 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=164 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=179 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=191 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=207 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=218 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=224 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=234 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=240 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=249 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=258 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=264 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=267 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=271 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=273 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=291 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=305 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=310 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=321 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=338 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=359 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=370 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=377 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=392 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=396 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=399 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=415 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=465 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=474 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=476 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=482 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=487 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=501 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=510 && yPixel<520) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=523 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=540 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=558 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=594 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=603 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=628 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=632 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=137 && xPixel<138 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=0 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=18 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=47 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=55 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=72 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=76 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=79 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=100 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=106 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=113 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=115 && yPixel<130) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=130 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=136 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=144 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=155 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=168 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=184 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=190 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=199 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=213 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=229 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=239 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=261 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=271 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=292 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=304 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=311 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=314 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=318 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=338 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=353 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=368 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=382 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=389 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=393 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=399 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=413 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=464 && yPixel<475) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=476 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=478 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=486 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=497 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=507 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=528 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=538 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=545 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=554 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=572 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=579 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=591 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=611 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=628 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=138 && xPixel<139 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=17 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=19 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=50 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=53 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=101 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=110 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=111 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=113 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=117 && yPixel<130) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=130 && yPixel<135) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=135 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=145 && yPixel<154) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=154 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=157 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=164 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=167 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=173 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=177 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=181 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=187 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=190 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=202 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=211 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=233 && yPixel<242) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=242 && yPixel<250) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=250 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=260 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=267 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=291 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=304 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=312 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=317 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=340 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=345 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=367 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=380 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=391 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=399 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=411 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=458 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=464 && yPixel<481) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=481 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=488 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=495 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=501 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=506 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=525 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=536 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=542 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=553 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=591 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=598 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=621 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=139 && xPixel<140 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=19 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=22 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=100 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=113 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=118 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=122 && yPixel<124) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=124 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=126 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=127 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=129 && yPixel<132) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=133 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=145 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=153 && yPixel<156) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=156 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=171 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=181 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=203 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=213 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=240 && yPixel<253) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=253 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=260 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=266 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=268 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=291 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=304 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=315 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=347 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=365 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=372 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=390 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=398 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=408 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=463 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=490 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=498 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=505 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=526 && yPixel<530) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=533 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=541 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=549 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=583 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=596 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=140 && xPixel<141 && yPixel>=620 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=22 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=27 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=52 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=101 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=123 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=145 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=151 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=160 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=170 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=177 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=206 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=215 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=236 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=256 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=261 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=267 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=291 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=297 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=312 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=316 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=346 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=363 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=370 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=385 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=398 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=406 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=456 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=463 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=483 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=500 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=504 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=521 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=529 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=540 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=544 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=564 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=597 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=608 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=619 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=141 && xPixel<142 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=0 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=23 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=28 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=80 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=104 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=118 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=120 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=122 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=124 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=151 && yPixel<156) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=156 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=201 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=220 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=224 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=237 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=256 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=290 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=295 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=298 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=307 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=315 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=346 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=362 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=369 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=381 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=397 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=404 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=455 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=463 && yPixel<478) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=478 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=493 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=499 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=516 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=523 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=526 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=543 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=564 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=580 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=595 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=616 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=142 && xPixel<143 && yPixel>=622 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=0 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=23 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=26 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=29 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=80 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=86 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=105 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=111 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=116 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=121 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=126 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=146 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=152 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=200 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=211 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=215 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=225 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=229 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=256 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=297 && yPixel<304) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=305 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=313 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=346 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=360 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=366 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=378 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=398 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=402 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=462 && yPixel<476) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=476 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=490 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=499 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=510 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=516 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=518 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=562 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=565 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=585 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=592 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=621 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=143 && xPixel<144 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=24 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=32 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=83 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=107 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=111 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=116 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=119 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=133 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=147 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=152 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=203 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=215 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=221 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=231 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=258 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=312 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=346 && yPixel<359) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=359 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=365 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=375 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=454 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=462 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=474 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=481 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=486 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=492 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=496 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=501 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=509 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=577 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=582 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=596 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=619 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=144 && xPixel<145 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=33 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=48 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=78 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=107 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=114 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=117 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=135 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=140 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=144 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=156 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=160 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=164 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=166 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=209 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=215 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=219 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=231 && yPixel<255) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=259 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=295 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=307 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=312 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=324 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=345 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=358 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=364 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=372 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=453 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=462 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=475 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=491 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=500 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=579 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=588 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=604 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=624 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=145 && xPixel<146 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=0 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=36 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=87 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=107 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=110 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=112 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=117 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=152 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=158 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=163 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=169 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=183 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=187 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=217 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=225 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=230 && yPixel<254) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=255 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=257 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=302 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=310 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=319 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=323 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=344 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=357 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=362 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=369 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=453 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=459 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=468 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=471 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=474 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=480 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=484 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=490 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=495 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=553 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=574 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=592 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=603 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=609 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=618 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=624 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=146 && xPixel<147 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=28 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=32 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=37 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=90 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=96 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=108 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=116 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=118 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=148 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=152 && yPixel<154) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=154 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=163 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=170 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=176 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=180 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=189 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=199 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=226 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=230 && yPixel<250) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=250 && yPixel<253) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=253 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=257 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=274 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=281 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=294 && yPixel<301) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=301 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=308 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=321 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=324 && yPixel<343) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=343 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=356 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=360 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=366 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=453 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=459 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=479 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=487 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=494 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=548 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=564 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=590 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=611 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=616 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=630 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=147 && xPixel<148 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=0 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=31 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=41 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=68 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=80 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=91 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=95 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=98 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=109 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=112 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=116 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=118 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=143 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=152 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=158 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=160 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=163 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=170 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=206 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=219 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=227 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=233 && yPixel<252) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=255 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=274 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=294 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=300 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=313 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=321 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=324 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=342 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=354 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=359 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=365 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=406 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=435 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=452 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=461 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=478 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=486 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=497 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=543 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=571 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=582 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=602 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=616 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=621 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=148 && xPixel<149 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=32 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=47 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=69 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=85 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=98 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=109 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=112 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=115 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=117 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=118 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=119 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=135 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=142 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=157 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=165 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=173 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=178 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=216 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=224 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=230 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=234 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=238 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=252 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=270 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=273 && yPixel<278) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=279 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=293 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=306 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=314 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=320 && yPixel<325) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=325 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=340 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=352 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=355 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=362 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=400 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=406 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=434 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=450 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=458 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=475 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=477 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=485 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=499 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=539 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=565 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=578 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=582 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=596 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=614 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=619 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=149 && xPixel<150 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=0 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=31 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=37 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=40 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=50 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=73 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=76 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=80 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=92 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=97 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=100 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=102 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=108 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=114 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=117 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=119 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=120 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=134 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=138 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=143 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=146 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=150 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=155 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=162 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=166 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=169 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=178 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=206 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=215 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=225 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=230 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=240 && yPixel<247) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=247 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=272 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=276 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=294 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=304 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=312 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=318 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=329 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=339 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=352 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=361 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=398 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=406 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=432 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=446 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=456 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=467 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=471 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=476 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=478 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=484 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=499 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=528 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=535 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=548 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=555 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=588 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=596 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=617 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=629 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=150 && xPixel<151 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=0 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=30 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=32 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=38 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=42 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=51 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=74 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=77 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=80 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=92 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=98 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=101 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=104 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=108 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=117 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=119 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=121 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=131 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=134 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=138 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=140 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=142 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=146 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=161 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=168 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=176 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=182 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=187 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=189 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=192 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=197 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=201 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=205 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=220 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=233 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=236 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=244 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=248 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=268 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=278 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=289 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=295 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=305 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=311 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=322 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=328 && yPixel<337) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=337 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=351 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=359 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=397 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=408 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=431 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=444 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=455 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=467 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=473 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=476 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=481 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=484 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=494 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=498 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=521 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=531 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=546 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=555 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=559 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=570 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=575 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=588 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=604 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=618 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=151 && xPixel<152 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=0 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=33 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=53 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=94 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=106 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=112 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=120 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=131 && yPixel<135) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=139 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=148 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=160 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=168 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=176 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=181 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=184 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=186 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=194 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=198 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=201 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=213 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=222 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=229 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=237 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=246 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=267 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=272 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=279 && yPixel<287) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=287 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=304 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=322 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=328 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=336 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=350 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=357 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=394 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=408 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=430 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=442 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=455 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=461 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=466 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=469 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=481 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=490 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=499 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=503 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=515 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=544 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=561 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=574 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=583 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=587 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=591 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=602 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=608 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=152 && xPixel<153 && yPixel>=618 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=32 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=53 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=95 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=107 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=120 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=124 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=137 && yPixel<138) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=138 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=147 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=161 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=164 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=168 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=174 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=179 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=190 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=194 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=200 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=218 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=223 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=227 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=231 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=237 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=247 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=267 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=270 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=278 && yPixel<283) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=283 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=289 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=295 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=303 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=312 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=323 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=327 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=333 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=348 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=355 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=392 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=406 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=429 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=442 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=450 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=458 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=461 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=466 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=468 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=480 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=499 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=502 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=517 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=533 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=578 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=587 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=612 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=618 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=153 && xPixel<154 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=0 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=31 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=51 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=53 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=57 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=64 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=71 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=94 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=99 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=107 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=128 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=146 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=160 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=173 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=182 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=194 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=198 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=203 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=211 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=219 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=228 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=237 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=249 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=264 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=267 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=288 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=295 && yPixel<301) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=307 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=314 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=321 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=330 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=344 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=346 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=352 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=392 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=404 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=422 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=425 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=440 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=450 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=454 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=460 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=470 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=483 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=496 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=500 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=514 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=526 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=568 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=581 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=589 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=621 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=154 && xPixel<155 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=0 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=40 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=43 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=45 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=62 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=65 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=100 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=108 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=110 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=111 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=124 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=130 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=134 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=138 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=153 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=168 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=174 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=182 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=186 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=197 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=206 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=219 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=230 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=250 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=262 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=265 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=276 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=295 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=301 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=313 && yPixel<322) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=322 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=345 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=350 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=391 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=402 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=424 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=438 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=451 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=453 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=461 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=470 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=481 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=492 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=499 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=515 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=524 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=535 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=552 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=567 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=581 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=592 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=607 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=155 && xPixel<156 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=0 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=33 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=38 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=42 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=54 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=58 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=64 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=66 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=67 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=69 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=98 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=103 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=108 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=114 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=117 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=124 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=142 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=145 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=151 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=169 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=177 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=186 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=213 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=218 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=225 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=233 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=251 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=262 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=264 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=274 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=311 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=321 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=343 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=347 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=390 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=401 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=434 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=460 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=469 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=482 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=494 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=501 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=508 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=519 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=524 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=527 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=545 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=571 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=578 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=603 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=616 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=624 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=156 && xPixel<157 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=0 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=35 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=37 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=39 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=42 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=45 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=54 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=58 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=61 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=64 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=71 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=114 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=117 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=124 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=141 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=152 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=169 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=175 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=186 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=190 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=222 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=232 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=250 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=262 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=264 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=273 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=298 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=321 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=345 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=389 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=400 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=432 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=465 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=470 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=472 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=478 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=483 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=519 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=556 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=568 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=584 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=601 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=619 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=629 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=157 && xPixel<158 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=0 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=40 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=56 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=62 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=65 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=69 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=73 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=115 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=119 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=122 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=126 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=144 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=152 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=169 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=171 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=175 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=184 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=187 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=189 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=206 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=211 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=220 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=233 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=245 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=260 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=264 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=272 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=291 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=297 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=320 && yPixel<338) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=340 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=342 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=381 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=387 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=400 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=431 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=460 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=469 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=475 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=483 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=522 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=526 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=561 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=568 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=575 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=581 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=602 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=610 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=617 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=622 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=158 && xPixel<159 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=0 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=43 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=65 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=73 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=102 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=117 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=120 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=123 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=125 && yPixel<127) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=128 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=139 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=148 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=153 && yPixel<156) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=158 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=164 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=171 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=176 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=186 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=211 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=216 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=219 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=225 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=244 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=262 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=264 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=270 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=278 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=280 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=294 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=321 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=341 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=385 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=398 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=414 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=418 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=429 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=466 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=468 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=481 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=532 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=554 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=577 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=597 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=604 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=629 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=159 && xPixel<160 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=0 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=44 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=46 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=59 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=66 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=72 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=74 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=105 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=120 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=135 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=139 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=143 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=146 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=155 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=167 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=173 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=179 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=182 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=184 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=209 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=219 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=244 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=263 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=269 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=275 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=280 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=293 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=319 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=337 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=340 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=385 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=393 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=408 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=413 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=418 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=428 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=448 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=466 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=489 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=517 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=520 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=529 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=550 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=558 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=572 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=597 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=608 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=618 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=160 && xPixel<161 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=0 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=46 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=60 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=64 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=74 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=101 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=105 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=131 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=134 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=140 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=142 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=146 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=152 && yPixel<154) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=154 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=167 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=176 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=183 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=203 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=223 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=234 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=244 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=263 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=268 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=272 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=281 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=284 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=290 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=317 && yPixel<332) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=332 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=338 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=381 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=392 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=412 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=417 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=426 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=448 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=464 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=487 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=493 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=517 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=523 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=556 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=566 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=578 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=612 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=623 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=161 && xPixel<162 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=0 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=47 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=60 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=63 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=75 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=105 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=120 && yPixel<132) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=133 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=169 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=176 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=183 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=203 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=216 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=230 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=236 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=244 && yPixel<259) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=259 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=262 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=272 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=275 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=316 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=337 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=385 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=404 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=415 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=424 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=454 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=491 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=500 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=506 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=518 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=536 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=542 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=551 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=560 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=571 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=594 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=609 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=162 && xPixel<163 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=0 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=47 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=61 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=64 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=69 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=72 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=76 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=118 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=145 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=151 && yPixel<154) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=154 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=169 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=179 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=183 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=207 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=214 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=221 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=232 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=236 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=243 && yPixel<259) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=259 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=262 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=269 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=316 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=336 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=389 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=403 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=414 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=424 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=446 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=450 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=489 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=497 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=508 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=519 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=537 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=542 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=551 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=561 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=571 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=582 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=593 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=603 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=163 && xPixel<164 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=0 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=49 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=64 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=70 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=77 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=117 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=143 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=169 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=180 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=188 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=195 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=209 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=218 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=221 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=227 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=236 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=245 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=263 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=267 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=270 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=313 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=334 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=387 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=400 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=412 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=421 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=447 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=450 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=497 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=507 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=517 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=537 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=542 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=549 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=573 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=581 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=593 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=603 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=628 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=632 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=164 && xPixel<165 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=0 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=50 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=68 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=71 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=77 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=113 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=115 && yPixel<131) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=131 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=136 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=140 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=149 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=165 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=169 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=175 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=180 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=189 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=191 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=195 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=207 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=217 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=226 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=234 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=246 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=257 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=265 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=271 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=276 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=304 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=310 && yPixel<325) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=327 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=333 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=354 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=365 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=386 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=399 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=410 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=418 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=503 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=505 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=513 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=537 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=545 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=570 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=585 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=603 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=624 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=630 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=165 && xPixel<166 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=0 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=50 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=54 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=58 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=63 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=72 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=76 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=78 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=80 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=107 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=126 && yPixel<128) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=130 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=134 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=137 && yPixel<138) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=138 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=145 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=151 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=155 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=161 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=170 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=174 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=205 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=217 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=220 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=225 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=233 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=247 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=257 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=263 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=269 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=275 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=303 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=311 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=323 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=326 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=331 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=349 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=355 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=362 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=364 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=381 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=384 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=390 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=396 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=408 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=419 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=510 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=537 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=554 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=561 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=572 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=589 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=629 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=166 && xPixel<167 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=0 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=51 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=57 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=61 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=66 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=69 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=72 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=78 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=83 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=106 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=125 && yPixel<132) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=132 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=143 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=160 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=202 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=207 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=216 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=219 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=228 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=235 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=238 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=247 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=258 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=268 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=275 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=297 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=317 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=324 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=330 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=348 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=354 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=358 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=366 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=378 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=381 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=390 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=396 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=407 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=419 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=433 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=510 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=547 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=556 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=561 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=570 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=586 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=601 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=614 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=620 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=167 && xPixel<168 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=0 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=48 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=51 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=53 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=58 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=65 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=68 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=74 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=76 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=81 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=95 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=122 && yPixel<125) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=125 && yPixel<129) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=129 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=138 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=143 && yPixel<154) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=154 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=161 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=183 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=189 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=192 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=197 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=201 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=208 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=228 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=232 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=237 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=247 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=258 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=272 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=302 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=304 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=310 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=321 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=328 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=337 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=345 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=358 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=361 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=365 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=394 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=406 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=417 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=434 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=509 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=539 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=548 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=555 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=574 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=587 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=604 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=168 && xPixel<169 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=0 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=49 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=51 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=58 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=69 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=71 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=76 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=80 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=101 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=125 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=127 && yPixel<129) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=129 && yPixel<132) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=134 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=140 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=144 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=147 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=161 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=181 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=188 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=208 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=217 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=229 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=237 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=247 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=258 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=270 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=276 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=285 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=304 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=312 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=318 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=325 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=339 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=344 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=354 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=362 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=386 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=394 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=404 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=416 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=451 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=505 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=555 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=570 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=575 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=583 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=601 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=620 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=629 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=169 && xPixel<170 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=0 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=51 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=59 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=66 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=67 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=69 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=82 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=87 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=99 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=102 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=129 && yPixel<135) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=135 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=144 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=148 && yPixel<156) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=156 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=161 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=168 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=178 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=186 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=197 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=215 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=225 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=229 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=235 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=246 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=256 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=275 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=302 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=317 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=323 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=339 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=343 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=359 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=383 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=395 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=403 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=417 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=449 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=451 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=500 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=541 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=553 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=569 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=581 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=627 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=170 && xPixel<171 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=0 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=82 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=86 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=90 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=93 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=101 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=131 && yPixel<134) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=134 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=137 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=143 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=155 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=161 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=168 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=181 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=184 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=187 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=195 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=207 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=215 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=227 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=234 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=247 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=257 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=270 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=275 && yPixel<282) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=302 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=322 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=335 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=341 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=358 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=371 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=378 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=395 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=400 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=413 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=417 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=423 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=428 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=503 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=542 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=552 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=569 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=580 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=589 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=592 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=598 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=619 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=171 && xPixel<172 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=0 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=87 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=90 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=93 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=102 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=105 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=136 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=151 && yPixel<154) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=154 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=156 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=160 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=182 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=187 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=195 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=208 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=224 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=228 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=234 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=245 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=249 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=256 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=281 && yPixel<286) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=299 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=302 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=306 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=311 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=321 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=329 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=340 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=361 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=368 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=382 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=398 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=410 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=418 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=501 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=537 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=542 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=558 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=566 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=582 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=611 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=172 && xPixel<173 && yPixel>=614 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=0 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=90 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=94 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=106 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=133 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=138 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=153 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=157 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=162 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=168 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=181 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=187 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=196 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=209 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=227 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=232 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=248 && yPixel<255) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=255 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=291 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=306 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=311 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=319 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=327 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=339 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=353 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=360 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=366 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=383 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=390 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=402 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=412 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=417 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=499 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=561 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=569 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=572 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=578 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=583 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=599 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=613 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=625 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=173 && xPixel<174 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=0 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=99 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=105 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=130 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b11000000,8'b11000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=152 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=155 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=165 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=179 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=191 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=198 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=206 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=232 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=250 && yPixel<254) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=254 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=297 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=306 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=311 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=317 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=326 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=339 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=351 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=358 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=361 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=364 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=388 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=398 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=416 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=423 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=497 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=546 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=553 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=570 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=576 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=615 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=622 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=629 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=174 && xPixel<175 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=0 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=99 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=105 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=109 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=124 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=130 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=143 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b11000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=151 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=158 && yPixel<160) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=160 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=163 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=175 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=178 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=187 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=200 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=234 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=252 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=294 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=299 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=306 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=310 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=316 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=323 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=339 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=343 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=349 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=361 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=378 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=383 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=384 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=395 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=411 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=421 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=494 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=525 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=530 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=535 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=558 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=570 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=577 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=586 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=596 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=616 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=620 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=628 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=175 && xPixel<176 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=0 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=106 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=109 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=123 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=137 && yPixel<142) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=144 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=148 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=159 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=187 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=195 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=198 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=234 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=251 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=284 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=294 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=301 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=307 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=321 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=331 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=354 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=359 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=394 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=406 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=420 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=425 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=491 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=529 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=531 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=554 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=564 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=574 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=604 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=625 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=176 && xPixel<177 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=0 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=100 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=107 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=109 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=110 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=111 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=123 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=137 && yPixel<143) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=143 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=162 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=174 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=183 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=187 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=198 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=237 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=252 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=277 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=299 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=305 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=319 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=331 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=343 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=357 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=376 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=386 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=396 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=402 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=408 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=420 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=432 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=461 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=487 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=517 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=529 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=535 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=543 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=546 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=577 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=592 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=596 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=611 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=177 && xPixel<178 && yPixel>=615 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=0 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=107 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=109 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=123 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=133 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=137 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=148 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=165 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=182 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=190 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=196 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=239 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=250 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=254 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=277 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=293 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=300 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=319 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=331 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=339 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=343 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=355 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=363 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=373 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=378 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=402 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=417 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=433 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=462 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=485 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=519 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=529 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=532 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=546 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=563 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=570 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=601 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=607 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=178 && xPixel<179 && yPixel>=619 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=0 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=102 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=108 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=121 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=124 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=130 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=147 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=166 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=175 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=181 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=190 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=199 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=239 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=244 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=250 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=254 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=278 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=282 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=297 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=301 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=308 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=319 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=327 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=335 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=342 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=354 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=361 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=367 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=369 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=373 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=398 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=407 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=416 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=426 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=432 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=461 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=484 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=544 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=550 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=564 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=570 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=586 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=590 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b11000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=609 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=617 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=633 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=179 && xPixel<180 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=0 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=102 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=106 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=121 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=126 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=130 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=167 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=177 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=181 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=185 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=190 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=195 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=239 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=241 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=245 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=252 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=260 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=278 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=305 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=317 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=327 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=342 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=354 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=359 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=362 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=373 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=406 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=415 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=420 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=424 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=432 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=439 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=445 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=449 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=462 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=483 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=520 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=534 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=544 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=553 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=568 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=582 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=586 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=601 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=609 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=180 && xPixel<181 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=0 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=100 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=106 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=112 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=121 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=126 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=130 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=166 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=182 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=189 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=195 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=245 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=252 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=261 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=277 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=297 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=315 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=323 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=344 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=360 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=395 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=413 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=417 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=421 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=428 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=432 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=439 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=459 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=479 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=517 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=533 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=544 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=548 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=552 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=567 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=579 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=583 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=600 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=605 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=624 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=181 && xPixel<182 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=0 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=101 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=111 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=121 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=124 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=127 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=129 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=165 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=175 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=181 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=244 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=251 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=256 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=262 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=270 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=277 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=296 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=312 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=321 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=336 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=340 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=383 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=392 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=397 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=404 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=415 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=421 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=427 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=437 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=451 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=459 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=471 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=517 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=529 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=542 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=551 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=556 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=567 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=581 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=602 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=621 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=182 && xPixel<183 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=0 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=101 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=110 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=165 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=181 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=243 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=248 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=251 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=259 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=262 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=270 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=277 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=281 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=288 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=295 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=309 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=321 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=338 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=361 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=365 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=376 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=380 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=390 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=396 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=405 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=416 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=422 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=429 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=436 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=450 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=467 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=500 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=508 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=518 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=524 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=541 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=579 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=597 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=615 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=620 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=183 && xPixel<184 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=0 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=98 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=109 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=160 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=176 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=179 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=225 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=235 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=241 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=248 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=258 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=264 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=269 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=277 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=281 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=293 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=298 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=304 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=308 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=317 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=332 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=361 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=368 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=375 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=380 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=391 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=401 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=422 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=460 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=494 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=508 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=518 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=520 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=536 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=549 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=553 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=561 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=582 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=184 && xPixel<185 && yPixel>=592 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=0 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=96 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=106 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=161 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=174 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=178 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=219 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=223 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=234 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=240 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=259 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=265 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=268 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=274 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=281 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=297 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=315 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=329 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=340 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=344 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=359 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=364 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=377 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=380 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=393 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=396 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=400 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=426 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=488 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=506 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=517 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=536 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=560 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=574 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=579 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=589 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=185 && xPixel<186 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=0 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=93 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=104 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=156 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=164 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=174 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=180 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=193 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=198 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=214 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=221 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=237 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=244 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=256 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=267 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=275 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=281 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=293 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=301 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=319 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=330 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=338 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=342 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=371 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=393 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=399 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=422 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=481 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=484 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=504 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=512 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=527 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=532 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=537 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=554 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=575 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=585 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=633 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=186 && xPixel<187 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=0 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=93 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=102 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=109 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=110 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=154 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=168 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=180 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=186 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=189 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=197 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=218 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=221 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=244 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=256 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=275 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=278 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=288 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=299 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=302 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=316 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=323 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=330 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=339 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=350 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=386 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=398 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=422 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=431 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=476 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=499 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=510 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=524 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=534 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=537 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=543 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=547 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=568 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=575 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=581 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=622 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=630 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=187 && xPixel<188 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=0 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=94 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=101 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=104 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=110 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=153 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=169 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=177 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=182 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=185 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=195 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=210 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=217 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=227 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=244 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=250 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=255 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=272 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=275 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=278 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=289 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=299 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=306 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=316 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=330 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=337 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=352 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=383 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=384 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=393 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=396 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=420 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=478 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=499 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=510 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=521 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=544 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=551 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=562 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=570 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=577 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=596 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=610 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=619 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=632 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=188 && xPixel<189 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=0 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=45 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=94 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=100 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=102 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=109 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=153 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=169 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=183 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=189 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=192 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=197 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=204 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=214 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=229 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=242 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=256 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=269 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=278 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=288 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=298 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=309 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=318 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=331 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=353 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=368 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=374 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=384 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=393 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=426 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=476 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=478 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=492 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=510 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=515 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=531 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=546 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=551 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=568 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=590 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=598 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=605 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=627 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=189 && xPixel<190 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=0 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=42 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=44 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=47 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=94 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=101 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=107 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=152 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=170 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=196 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=205 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=212 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=231 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=239 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=256 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=269 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=278 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=291 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=298 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=304 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=307 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=318 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=331 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=350 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=368 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=379 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=386 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=390 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=419 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=423 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=428 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=477 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=493 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=511 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=529 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=542 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=550 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=557 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=564 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=586 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=591 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=601 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=623 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=631 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=190 && xPixel<191 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=0 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=41 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=43 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=50 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=95 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=101 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=107 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=153 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=171 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=176 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=183 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=193 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=197 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=205 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=210 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=219 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=237 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=256 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=268 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=278 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=288 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=301 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=307 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=317 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=354 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=380 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=386 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=436 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=490 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=504 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=522 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=533 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=549 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=573 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=580 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=586 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=591 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=597 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=191 && xPixel<192 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=0 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=40 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=42 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=53 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=94 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=101 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=107 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=150 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=176 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=183 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=193 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=198 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=200 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=208 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=215 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=231 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=235 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=242 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=288 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=302 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=320 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=336 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=383 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=437 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=500 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=517 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=528 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=533 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=538 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=549 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=566 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=583 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=589 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=595 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=615 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=627 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=192 && xPixel<193 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=0 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=41 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=55 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=94 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=102 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=107 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=148 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=172 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=179 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=184 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=189 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=192 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=200 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=207 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=212 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=231 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=236 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=244 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=268 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=288 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=292 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=300 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=309 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=321 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=374 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=437 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=440 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=443 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=447 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=450 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=499 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=514 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=523 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=535 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=541 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=549 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=576 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=586 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=602 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=608 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=622 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=193 && xPixel<194 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=0 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=41 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=56 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=93 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=102 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=111 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=148 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=178 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=183 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=191 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=199 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=209 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=235 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=255 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=262 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=284 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=291 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=304 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=309 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=322 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=373 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=437 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=444 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=447 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=456 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=499 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=512 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=524 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=529 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=540 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=548 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=602 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=606 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=618 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=194 && xPixel<195 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=5 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=10 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=41 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=58 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=93 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=102 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=116 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=148 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=177 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=182 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=186 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=213 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=236 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=257 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=261 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=280 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=283 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=290 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=305 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=309 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=348 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=372 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=437 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=442 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=449 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=455 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=497 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=515 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=522 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=531 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=539 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=545 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=559 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=563 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=576 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=586 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=599 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=611 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=621 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=634 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=195 && xPixel<196 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=3 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=5 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=7 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=17 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=19 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=41 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=60 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=92 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=102 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=120 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=148 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=176 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=179 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=186 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=196 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=205 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=213 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=280 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=283 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=287 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=290 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=309 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=317 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=438 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=446 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=452 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=461 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=495 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=511 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=527 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=533 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=542 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=553 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=565 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=573 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=594 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=602 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=620 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=196 && xPixel<197 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=5 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=15 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=19 && yPixel<22) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=22 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=40 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=42 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=59 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=65 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=91 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=103 && yPixel<127) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=127 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=149 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=178 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=182 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=185 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=193 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=196 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=211 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=217 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=282 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=299 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=309 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=317 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=356 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=361 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=431 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=441 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=451 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=461 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=481 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=492 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=508 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=530 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=551 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=563 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=568 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=582 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=589 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=591 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=606 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=619 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=627 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=197 && xPixel<198 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=3 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=8 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=23 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=26 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=43 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=61 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=64 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=66 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=88 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=98 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=101 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=107 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=118 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=119 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=148 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=181 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=192 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=197 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=210 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=216 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=245 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=265 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=267 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=270 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=288 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=294 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=301 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=305 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=313 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=341 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=351 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=359 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=435 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=453 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=462 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=466 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=471 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=484 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=505 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=527 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=531 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=546 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=577 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=582 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=587 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=608 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=617 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=620 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=198 && xPixel<199 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=2 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=3 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=8 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=26 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=33 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=38 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=47 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=68 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=87 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=98 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=107 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=125 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=133 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=148 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=180 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=192 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=196 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=206 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=216 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=221 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=252 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=264 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=276 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=288 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=292 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=304 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=319 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=329 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=345 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=355 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=467 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=472 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=478 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=499 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=526 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=541 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=568 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=573 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=583 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=593 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=607 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=618 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=627 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=199 && xPixel<200 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=6 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=29 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=47 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=70 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=74 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=86 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=101 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=108 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=116 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=117 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=123 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=128 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=131 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=150 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=178 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=193 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=226 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=248 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=257 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=264 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=272 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=276 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=284 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=291 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=307 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=319 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=329 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=490 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=517 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=528 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=540 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=577 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=599 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=605 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=612 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=621 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=630 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=200 && xPixel<201 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=2 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=31 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=34 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=47 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=73 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=77 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=83 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=98 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=103 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=109 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=123 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=128 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=136 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=149 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=172 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=177 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=220 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=229 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=241 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=244 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=247 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=258 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=264 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=270 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=276 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=287 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=302 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=306 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=319 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=329 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=467 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=486 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=536 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=557 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=568 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=576 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=600 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=613 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=201 && xPixel<202 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=3 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=33 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=51 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=72 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=98 && yPixel<104) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=104 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=110 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=120 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=124 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=138 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=148 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=169 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=173 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=176 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=217 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=222 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=233 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=241 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=257 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=264 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=269 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=280 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=295 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=306 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=328 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=482 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=527 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=534 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=546 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=550 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=554 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=565 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=575 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=582 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=587 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=593 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=610 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=615 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=620 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=202 && xPixel<203 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=3 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=33 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=49 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=72 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=98 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=105 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=112 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=123 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=173 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=205 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=216 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=222 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=234 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=247 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=261 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=269 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=281 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=287 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=297 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=305 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=320 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=329 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=351 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=481 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=520 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=526 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=530 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=548 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=564 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=571 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=576 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=592 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=602 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=606 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=616 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=632 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=203 && xPixel<204 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=5 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=32 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=36 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=52 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=57 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=61 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=73 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=75 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=96 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=106 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=114 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=124 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=135 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=144 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=150 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=171 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=174 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=202 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=221 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=238 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=248 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=253 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=261 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=268 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=272 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=285 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=292 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=302 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=320 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=326 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=352 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=477 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=514 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=522 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=536 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=544 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=560 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=576 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=587 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=591 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=602 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=617 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=622 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=204 && xPixel<205 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=4 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=34 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=52 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=56 && yPixel<60) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=60 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=64 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=74 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=77 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=96 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=106 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=116 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=125 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=131 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=137 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=139 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=174 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=200 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=216 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=222 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=242 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=249 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=253 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=265 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=272 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=285 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=291 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=295 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=317 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=323 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=350 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=356 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=472 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=510 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=518 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=542 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=547 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=552 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=569 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=591 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=598 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=613 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=620 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=630 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=205 && xPixel<206 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=4 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=36 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=52 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=59 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=65 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=72 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=77 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=98 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=107 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=117 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=121 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=123 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=129 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=153 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=178 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=200 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=214 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=219 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=222 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=246 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=249 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=264 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=271 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=285 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=290 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=322 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=342 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=469 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=499 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=510 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=525 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=547 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=551 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=569 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=573 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=578 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=585 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=589 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=610 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=615 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=206 && xPixel<207 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=10 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=39 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=52 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=55 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=69 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=74 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=77 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=94 && yPixel<97) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=99 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=108 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=117 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=121 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=129 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=155 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=173 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=179 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=199 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=213 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=231 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=246 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=252 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=278 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=285 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=294 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=322 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=361 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=466 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=496 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=511 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=523 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=535 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=546 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=565 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=578 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=585 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=608 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=623 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=207 && xPixel<208 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=12 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=40 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=52 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=54 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=74 && yPixel<77) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=77 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=82 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=94 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=99 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=109 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=118 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=126 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=145 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=149 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=157 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=173 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=180 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=199 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=213 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=229 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=244 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=259 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=265 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=272 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=284 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=289 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=300 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=310 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=321 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=353 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=366 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=403 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=463 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=492 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=497 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=511 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=526 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=550 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=563 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=570 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=582 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=608 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=620 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=208 && xPixel<209 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=18 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=45 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=55 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=61 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=66 && yPixel<78) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=78 && yPixel<86) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=86 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=91 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=95 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=99 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=111 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=119 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=124 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=152 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=168 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=173 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=180 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=198 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=211 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=220 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=224 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=231 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=241 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=247 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=253 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=261 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=267 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=269 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=284 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=298 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=307 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=342 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=353 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=363 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=461 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=495 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=509 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=532 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=542 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=551 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=560 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=564 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=574 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=577 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=593 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=612 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=619 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=629 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=632 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=209 && xPixel<210 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=14 && yPixel<16) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=17 && yPixel<20) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=23 && yPixel<29) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=29 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=46 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=53 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=56 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=59 && yPixel<71) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=71 && yPixel<83) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=85 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=91 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=95 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=98 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=112 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=119 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=126 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=128 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=166 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=169 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=172 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=180 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=198 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=210 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=215 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=238 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=247 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=261 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=266 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=282 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=287 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=290 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=301 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=312 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=324 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=335 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=344 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=407 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=459 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=486 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=495 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=500 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=527 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=553 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=559 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b11000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=571 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=581 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=587 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=619 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=627 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=210 && xPixel<211 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=9 && yPixel<24) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=26 && yPixel<32) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=32 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=46 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=52 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=56 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=59 && yPixel<75) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=75 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=90 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=98 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=114 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=119 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=122 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=131 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=165 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=176 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=180 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=196 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=209 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=217 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=241 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=267 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=271 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=275 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=289 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=300 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=311 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=323 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=331 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=341 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=457 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=484 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=491 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=495 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=498 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=507 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=529 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=556 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=565 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=583 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=603 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=617 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=211 && xPixel<212 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=9 && yPixel<26) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=30 && yPixel<37) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=37 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=42 && yPixel<45) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=45 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=56 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=59 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=73 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=98 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=115 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=120 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=124 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=127 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=132 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=162 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=165 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=176 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=181 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=194 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=210 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=218 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=226 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=244 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=255 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=265 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=289 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=306 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=313 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=319 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=323 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=332 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=337 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=347 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=352 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=457 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=480 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=491 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=497 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=502 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=506 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=517 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b11000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=557 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=562 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=578 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=588 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=603 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=611 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=212 && xPixel<213 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=11 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=34 && yPixel<47) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=47 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=56 && yPixel<60) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=60 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=73 && yPixel<88) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=88 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=95 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=98 && yPixel<116) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=116 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=120 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=124 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=126 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=130 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=137 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=163 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=176 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=181 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=194 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=208 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=218 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=226 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=246 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=259 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=274 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=294 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=306 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=318 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=336 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=341 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=351 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=457 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=477 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=489 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=496 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=512 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=527 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=548 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=558 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=574 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=580 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=597 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=606 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=617 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=213 && xPixel<214 && yPixel>=620 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=12 && yPixel<33) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=33 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=49 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=55 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=61 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=73 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=79 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=82 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=85 && yPixel<90) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=90 && yPixel<117) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=117 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=121 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=124 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=126 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=129 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=143 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=153 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=163 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=175 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=183 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=194 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=207 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=230 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=249 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=256 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=262 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=277 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=300 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=313 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=331 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=457 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=474 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=479 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=504 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=506 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=513 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=543 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=545 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=555 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=570 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=575 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=601 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=616 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=214 && xPixel<215 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=13 && yPixel<32) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=32 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=55 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=62 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=74 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=79 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=82 && yPixel<86) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=86 && yPixel<89) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=89 && yPixel<93) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=93 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=118 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=121 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=126 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=136 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=153 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=158 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=175 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=184 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=194 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=206 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=221 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=230 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=261 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=275 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=292 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=299 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=458 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=471 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=479 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=493 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=512 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=535 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=542 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=551 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=566 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=572 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=603 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=610 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=626 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=215 && xPixel<216 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=0 && yPixel<15) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=15 && yPixel<32) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=34 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=62 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=74 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=82 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=84 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=87 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=91 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=96 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=118 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=122 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=130 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=133 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=144 && yPixel<148) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=148 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=152 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=157 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=173 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=185 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=193 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=204 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=213 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=224 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=254 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=310 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=468 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=489 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=496 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=499 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=503 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=518 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=532 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=539 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=549 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=569 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=591 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=600 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=603 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=614 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=617 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=216 && xPixel<217 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=0 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=16 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=34 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=62 && yPixel<75) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=75 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=79 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=84 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=93 && yPixel<97) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=97 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=119 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=122 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=133 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=147 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=166 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=191 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=205 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=209 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=225 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=251 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=266 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=273 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=279 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=295 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=298 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=331 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=469 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=484 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=498 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=502 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=533 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=548 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=560 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=566 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=597 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=603 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=610 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=625 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=217 && xPixel<218 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=3 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=18 && yPixel<32) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=32 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=57 && yPixel<63) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=63 && yPixel<75) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=75 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=84 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=98 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=119 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=122 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=146 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=165 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=208 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=224 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=241 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=245 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=252 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=267 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=273 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=278 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=286 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=294 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=322 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=472 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=487 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=491 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=502 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=505 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=518 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=520 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=524 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=530 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=535 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=546 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=555 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=562 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=580 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=587 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=597 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=609 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=622 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=630 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=218 && xPixel<219 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=6 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=18 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=34 && yPixel<63) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=63 && yPixel<75) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=75 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=84 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=98 && yPixel<100) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=100 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=118 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=122 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=147 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=164 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=202 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=208 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=211 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=218 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=224 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=242 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=254 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=263 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=273 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=288 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=294 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=315 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=322 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=327 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=366 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=466 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=482 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=485 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=493 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=502 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=513 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=525 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=530 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=538 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=549 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=559 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=574 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=581 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=587 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=601 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=616 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=626 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=219 && xPixel<220 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=8 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=20 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=34 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=64 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=74 && yPixel<84) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=84 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=98 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=101 && yPixel<118) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=118 && yPixel<122) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=122 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=153 && yPixel<164) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=164 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=201 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=211 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=216 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=219 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=225 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=231 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=241 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=252 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=255 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=262 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=265 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=269 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=289 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=305 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=336 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=365 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=463 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=482 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=485 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=491 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=500 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=504 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=509 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=516 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=526 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=547 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=558 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=576 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=585 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=595 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=612 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b10000000};
	if(xPixel>=220 && xPixel<221 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=10 && yPixel<21) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=21 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=34 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=65 && yPixel<73) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=73 && yPixel<82) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=82 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=100 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=103 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=115 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=121 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=157 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=165 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=200 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=211 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=219 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=227 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=231 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=266 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=279 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=284 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=292 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=325 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=328 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=353 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=356 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=362 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=370 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=460 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=481 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=491 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=497 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=505 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=509 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=521 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=530 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=544 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=547 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=556 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=566 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=580 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=590 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=604 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=612 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=221 && xPixel<222 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=12 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=23 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=34 && yPixel<36) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=37 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=66 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=72 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=81 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=102 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=106 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=121 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=154 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=158 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=167 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=200 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=210 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=215 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=219 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=223 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=226 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=229 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=254 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=267 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=279 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=291 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=306 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=313 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=318 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=329 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=347 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=363 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=368 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=371 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=373 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=383 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=458 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=478 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=483 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=491 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=499 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=517 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=525 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=530 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=534 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=539 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=558 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=575 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=580 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=592 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=601 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=607 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=619 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=222 && xPixel<223 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=13 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=25 && yPixel<34) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=34 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=68 && yPixel<71) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=71 && yPixel<78) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=78 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=104 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=109 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=115 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=120 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=161 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=168 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=208 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=222 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=228 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=244 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=251 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=255 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=259 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=279 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=303 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=308 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=322 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=335 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=345 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=356 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=366 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=370 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=385 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=454 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=484 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=489 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=513 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=523 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=531 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=534 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=544 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=550 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=580 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=588 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=595 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=602 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=613 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=623 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=223 && xPixel<224 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=0 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=15 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=26 && yPixel<36) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=36 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=55 && yPixel<60) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=62 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=65 && yPixel<67) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=67 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=72 && yPixel<78) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=78 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=107 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=112 && yPixel<115) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=115 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=119 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=152 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=155 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=162 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=169 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=206 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=219 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=248 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=271 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=286 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=296 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=307 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=319 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=327 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=343 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=362 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=367 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=383 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=402 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=451 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=476 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=485 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=499 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=503 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=515 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=518 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=528 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=542 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=560 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=574 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=590 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=595 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b11000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=608 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=613 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=224 && xPixel<225 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=17 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=28 && yPixel<38) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=38 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=53 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=61 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=65 && yPixel<67) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=70 && yPixel<79) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=79 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=110 && yPixel<119) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=119 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=161 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=170 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=206 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=216 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=246 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=253 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=265 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=283 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=290 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=301 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=331 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=342 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=359 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=366 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=370 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=379 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=385 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=394 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=401 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=449 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=475 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=479 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=486 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=499 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=514 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=531 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=554 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=588 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=603 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=609 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=614 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=619 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=625 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=225 && xPixel<226 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=19 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=30 && yPixel<38) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=38 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=54 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=58 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=64 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=66 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=72 && yPixel<80) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=80 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=113 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=120 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=155 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=162 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=171 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=183 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=206 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=217 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=220 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=246 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=259 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=267 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=273 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=300 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=308 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=326 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=336 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=349 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=358 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=365 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=395 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=446 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=472 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=474 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=477 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=496 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=503 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=507 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=516 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=547 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=558 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=577 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=584 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=597 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=226 && xPixel<227 && yPixel>=610 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=22 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=32 && yPixel<40) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=40 && yPixel<52) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=52 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=57 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=62 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=65 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=72 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=77 && yPixel<81) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=81 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=117 && yPixel<120) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=120 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=156 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=164 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=171 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=181 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=184 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=191 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=197 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=206 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=223 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=258 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=266 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=268 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=276 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=280 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=318 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=353 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=361 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=409 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=443 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=470 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=472 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=480 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=490 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=500 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=506 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=519 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=523 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=540 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=550 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=555 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=578 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=592 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=608 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=227 && xPixel<228 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=24 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=34 && yPixel<40) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=40 && yPixel<52) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=52 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=61 && yPixel<63) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=63 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=69 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=168 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=173 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=180 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=191 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=206 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=222 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=256 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=266 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=268 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=272 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=283 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=285 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=303 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=322 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=328 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=359 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=362 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=365 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=375 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=384 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=391 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=397 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=409 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=440 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=467 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=472 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=482 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=488 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=493 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=497 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=501 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=505 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=514 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=533 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=540 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=550 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=574 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=584 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=589 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=601 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=609 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=228 && xPixel<229 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=0 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=25 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=35 && yPixel<41) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=41 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=53 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=68 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=171 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=176 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=179 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=191 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=207 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=223 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=255 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=267 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=301 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=308 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=314 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=321 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=328 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=351 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=355 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=359 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=362 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=366 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=415 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=437 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=458 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=462 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=470 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=472 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=481 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=486 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=496 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=501 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=519 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=531 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=546 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=555 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=564 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=577 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=597 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=229 && xPixel<230 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=26 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=33 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=36 && yPixel<42) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=42 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=55 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=173 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=191 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=207 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=224 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=254 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=268 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=274 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=281 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=315 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=326 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=344 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=353 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=423 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=435 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=459 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=464 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=472 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=477 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=479 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=487 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=495 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=506 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=516 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=525 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=534 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=542 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=559 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=577 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=589 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=604 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=610 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=230 && xPixel<231 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=26 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=32 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=36 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=43 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=57 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=166 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=175 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=186 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=191 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=203 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=208 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=224 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=254 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=266 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=271 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=286 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=309 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=314 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=325 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=338 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=421 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=433 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=457 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=460 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=473 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=477 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=488 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=500 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=508 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=514 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=527 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=529 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=537 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=549 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=571 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=576 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=599 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=619 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=627 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=231 && xPixel<232 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=26 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=33 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=36 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=43 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=50 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=58 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=176 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=191 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=203 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=208 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=224 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=254 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=265 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=267 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=286 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=300 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=321 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=329 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=358 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=370 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=419 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=432 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=454 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=458 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=471 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=477 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=483 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=499 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=511 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=523 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=530 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=580 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=593 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=608 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=617 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=232 && xPixel<233 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=24 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=28 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=32 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=35 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=37 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=43 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=49 && yPixel<51) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=51 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=61 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=177 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=223 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=252 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=260 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=265 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=267 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=273 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=279 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=283 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=293 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=315 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=328 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=346 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=360 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=364 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=422 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=432 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=449 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=453 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=459 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=472 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=505 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=536 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=550 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=556 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=564 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=608 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=624 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=233 && xPixel<234 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=24 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=28 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=34 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=38 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=43 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=49 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=53 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=64 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=178 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=222 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=252 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=259 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=267 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=271 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=279 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=284 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=300 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=311 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=325 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=343 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=348 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=430 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=447 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=451 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=454 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=467 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=505 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=529 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=538 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=545 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=569 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=582 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=586 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=601 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=620 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=234 && xPixel<235 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=26 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=43 && yPixel<50) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=50 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=54 && yPixel<67) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=67 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=163 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=183 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=188 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=223 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=252 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=261 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=281 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=292 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=304 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=320 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=343 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=445 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=448 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=464 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=496 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=522 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=530 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=534 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=539 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=549 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=573 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=582 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=592 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=611 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=235 && xPixel<236 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=0 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=26 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=40 && yPixel<45) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=45 && yPixel<51) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=51 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=53 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=55 && yPixel<69) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=69 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=169 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=179 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=190 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=223 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=249 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=260 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=281 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=298 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=306 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=319 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=337 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=444 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=448 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=452 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=458 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=481 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=489 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=495 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=513 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=515 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=530 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=537 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=553 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=559 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=568 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=580 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=588 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=597 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=619 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=236 && xPixel<237 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=27 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=42 && yPixel<49) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=49 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=68 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=159 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=169 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=193 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=223 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=249 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=255 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=258 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=279 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=298 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=307 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=318 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=322 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=329 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=339 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=451 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=455 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=464 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=474 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=490 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=522 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=526 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=534 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=543 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=552 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=558 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=566 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=583 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=602 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=619 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=634 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=237 && xPixel<238 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=0 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=30 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=44 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=53 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=66 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=169 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=196 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=223 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=253 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=269 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=293 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=309 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=314 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=320 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=324 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=350 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=376 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=436 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=443 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=449 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=462 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=468 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=471 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=519 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=537 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=548 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=573 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=607 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=617 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=629 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=238 && xPixel<239 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=32 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=46 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=54 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=66 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=150 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=158 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=161 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=164 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=168 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=176 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=190 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=195 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=223 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=252 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=268 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=298 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=305 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=311 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=338 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=344 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=351 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=394 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=401 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=434 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=444 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=447 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=457 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=466 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=502 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=505 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=514 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=535 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=563 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=601 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=618 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=239 && xPixel<240 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=0 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=34 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=48 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=56 && yPixel<67) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=67 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=151 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=165 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=170 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=196 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=223 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=233 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=236 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=252 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=271 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=277 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=281 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=302 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=311 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=340 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=349 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=363 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=384 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=391 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=398 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=430 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=443 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=458 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=466 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=471 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=474 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=523 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=545 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=561 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=579 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=601 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=240 && xPixel<241 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=0 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=36 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=50 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=58 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=68 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=151 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=160 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=162 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=196 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=225 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=239 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=252 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=283 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=298 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=311 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=337 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=359 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=384 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=385 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=392 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=404 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=412 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=421 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=439 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=447 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=451 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=457 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=466 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=472 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=477 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=488 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=496 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=517 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=546 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=555 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=560 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=564 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=572 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=588 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=591 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=614 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=623 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=241 && xPixel<242 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=0 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=38 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=50 && yPixel<53) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=53 && yPixel<54) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=58 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=70 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=144 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=164 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=186 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=196 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=217 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=241 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=252 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=282 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=290 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=304 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=337 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=388 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=393 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=403 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=408 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=412 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=419 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=432 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=447 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=456 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=460 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=464 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=501 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=504 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=509 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=513 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=516 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=521 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=531 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=538 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=550 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=562 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=590 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=594 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=613 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=242 && xPixel<243 && yPixel>=626 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=0 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=41 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=51 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=58 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=70 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=144 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=163 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=195 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=217 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=243 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=252 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=285 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=300 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=319 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=327 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=331 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=348 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=359 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=381 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=394 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=401 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=413 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=416 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=425 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=447 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b11000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=460 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=472 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=474 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=484 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=499 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=512 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=525 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=542 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=547 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=566 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=592 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=609 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=622 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=243 && xPixel<244 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=0 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=34 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=45 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=61 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=64 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=68 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=165 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=177 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=182 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=190 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=203 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=217 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=242 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=252 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=256 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=282 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=297 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=318 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=338 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=348 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=361 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=379 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=383 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=388 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=405 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=411 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=416 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=441 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=446 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=457 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=473 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=509 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=512 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=519 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=527 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=539 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=546 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=563 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=595 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=601 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=619 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=626 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=244 && xPixel<245 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=0 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=35 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=47 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=165 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=182 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=190 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=203 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=217 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=241 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=256 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=299 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=308 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=314 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=334 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=380 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=386 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=393 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=398 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=410 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=415 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=432 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=438 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=444 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=505 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=515 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=524 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=530 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=542 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=564 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=597 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=245 && xPixel<246 && yPixel>=611 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=32 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=39 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=52 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=165 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=183 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=190 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=217 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=239 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=251 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=255 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=310 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=320 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=329 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=336 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=342 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=346 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=354 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=371 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=375 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=380 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=384 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=389 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=403 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=410 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=436 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=457 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=494 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=498 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=504 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=511 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=522 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=533 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=536 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=548 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=566 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=588 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=595 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=620 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=246 && xPixel<247 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=0 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=33 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=38 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=50 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=53 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=56 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=60 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=63 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=67 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=82 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=84 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=87 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=163 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=167 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=174 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=183 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=216 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=227 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=238 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=254 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=313 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=340 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=350 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=379 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=385 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=388 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=425 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=432 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=442 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=447 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=497 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=530 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=537 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=545 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=554 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=574 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=580 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=593 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=605 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=616 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=247 && xPixel<248 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=0 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=35 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=41 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=44 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=61 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=65 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=71 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=77 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=88 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=162 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=172 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=183 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=186 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=223 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=226 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=232 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=238 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=252 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=311 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=314 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=318 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=325 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=336 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=342 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=370 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=386 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=408 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b11000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=441 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=493 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=520 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=526 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=533 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=546 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=556 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=567 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=578 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=600 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=619 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=625 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=629 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=633 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=248 && xPixel<249 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=0 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=35 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=57 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=71 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=78 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=89 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=162 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=186 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=206 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=220 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=225 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=233 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=238 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=250 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=315 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=325 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=334 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=340 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=363 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=373 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=394 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=407 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=425 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=438 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=481 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=483 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=509 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=514 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=532 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=534 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=539 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=554 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=567 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=598 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=604 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=609 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=618 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=624 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=249 && xPixel<250 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=0 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=36 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=73 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=78 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=90 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=163 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=183 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=185 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=213 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=229 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=234 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=242 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=249 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=317 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=322 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=329 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=339 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=346 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=362 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=365 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=367 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=369 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=377 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=400 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=414 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=426 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=470 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=494 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=503 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=525 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=533 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=571 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=579 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=586 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=597 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=616 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=624 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=250 && xPixel<251 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=0 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=36 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=76 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=92 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=165 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=170 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=173 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=181 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=211 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=226 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=233 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=245 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=252 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=281 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=284 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=314 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=325 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=328 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=334 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=345 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=353 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=358 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=372 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=391 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=399 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=407 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=412 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b11000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=418 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=426 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=462 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=474 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=484 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=495 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=521 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=526 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=530 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=547 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=558 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=571 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=589 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=616 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=251 && xPixel<252 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=0 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=37 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=95 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=123 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=166 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=169 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=176 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=182 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=211 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=226 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=241 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=247 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=250 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=255 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=260 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=267 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=273 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=276 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=281 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=318 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=331 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=354 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=380 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=384 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=401 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=405 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=409 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b11000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=418 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=440 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=456 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=470 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=474 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=492 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=516 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=536 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=556 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=616 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=252 && xPixel<253 && yPixel>=621 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=0 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=39 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=93 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=122 && yPixel<126) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=126 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=165 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=169 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=176 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=183 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=211 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=225 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=240 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=260 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=265 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=274 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=280 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=310 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=318 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=324 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=384 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=392 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=404 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=462 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=480 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=486 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=497 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=509 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=524 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=529 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=532 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=543 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=554 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=615 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=626 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=253 && xPixel<254 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=0 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=41 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=91 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=122 && yPixel<128) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=128 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=170 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=173 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=177 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=184 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=211 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=224 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=239 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=271 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=274 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=279 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=292 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=306 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=311 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=323 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=326 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=459 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=464 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=472 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=474 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=484 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=486 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=494 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=498 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=502 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=512 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=517 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=526 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=544 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=609 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=254 && xPixel<255 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=0 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=40 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=43 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=80 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=91 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=125 && yPixel<131) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=131 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=150 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=169 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=181 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=213 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=221 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=238 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=260 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=265 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=269 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=274 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=278 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=290 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=294 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=311 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=324 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=391 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=398 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=461 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=465 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=478 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=491 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=494 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=500 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=508 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=514 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=517 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=522 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=547 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=559 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=611 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=616 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=621 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=255 && xPixel<256 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=0 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=41 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=44 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=80 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=87 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=88 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=96 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=152 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=178 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=191 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=193 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=228 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=255 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=267 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=270 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=273 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=277 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=288 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=310 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=313 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=327 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=382 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=389 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=394 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=397 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=405 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=458 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=462 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=466 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=469 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=482 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=510 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=537 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=541 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=556 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=597 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=607 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=611 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=256 && xPixel<257 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=13 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=16 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=20 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=43 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=47 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=65 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=82 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=84 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=86 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=97 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=177 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=225 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=241 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=254 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=264 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=277 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=286 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=296 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=324 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=407 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=410 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=453 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=463 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=467 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=480 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=511 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=537 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=554 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=567 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=588 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=610 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=257 && xPixel<258 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=13 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=18 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=26 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=45 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=49 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=97 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=166 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=172 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=176 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=196 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=208 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=219 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=233 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=237 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=243 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=248 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=264 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=267 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=272 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=288 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=318 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=336 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=381 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=384 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=397 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=418 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=457 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=462 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=479 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=498 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=500 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=507 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=517 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=523 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=528 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=535 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=544 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=549 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=567 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=577 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=586 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=258 && xPixel<259 && yPixel>=610 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=17 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=22 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=24 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=29 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=47 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=90 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=95 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=166 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=176 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=195 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=208 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=220 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=233 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=247 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=274 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=278 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=288 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=311 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=320 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=334 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=347 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=351 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=360 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=364 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=394 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=405 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=410 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=418 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=421 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=447 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=449 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=451 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=466 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=472 && yPixel<477) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=477 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=484 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=506 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=523 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=530 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=550 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=552 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=577 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=587 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=596 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=607 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=259 && xPixel<260 && yPixel>=623 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=20 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=25 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=30 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=36 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=52 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=89 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=94 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=164 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=173 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=178 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=185 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=192 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=215 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=274 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=279 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=293 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=317 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=323 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=334 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=338 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=354 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=357 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=362 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=374 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=384 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=391 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=402 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=417 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=431 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=433 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=440 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=444 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=464 && yPixel<468) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=468 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=469 && yPixel<482) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=482 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=490 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=497 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=504 && yPixel<519) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=519 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=530 && yPixel<532) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=533 && yPixel<545) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=571 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=580 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=588 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=619 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=260 && xPixel<261 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=22 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=37 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=58 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=62 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=64 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=96 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=166 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=173 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=217 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=240 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=272 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=293 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=304 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=315 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=329 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=344 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=348 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=354 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=360 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=378 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=389 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=411 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=422 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=433 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=443 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=450 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=462 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=491 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=504 && yPixel<523) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=527 && yPixel<546) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=558 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=574 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=588 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=261 && xPixel<262 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=18 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=47 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=51 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=71 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=102 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=214 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=220 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=229 && yPixel<245) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=245 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=277 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=286 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=300 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=304 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=311 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=320 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=328 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=333 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=344 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=355 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=373 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=375 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=378 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=391 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=416 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=427 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=438 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=460 && yPixel<464) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=465 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=497 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=500 && yPixel<525) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=526 && yPixel<546) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=616 && yPixel<628) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=262 && xPixel<263 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=15 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=19 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=75 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=107 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=214 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=228 && yPixel<254) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=255 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=257 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=271 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=281 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=284 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=310 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=317 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=327 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=333 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=355 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=388 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=395 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=408 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=411 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=435 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=458 && yPixel<464) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=465 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=496 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=499 && yPixel<551) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=565 && yPixel<570) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=584 && yPixel<588) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=603 && yPixel<632) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=263 && xPixel<264 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=12 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=26 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=78 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=82 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=115 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=260 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=275 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=283 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=302 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=308 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=320 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=327 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=341 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=346 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=360 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=395 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=407 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=435 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=457 && yPixel<463) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=464 && yPixel<493) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=497 && yPixel<506) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=507 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=516 && yPixel<538) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=539 && yPixel<555) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=565 && yPixel<572) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=582 && yPixel<594) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=264 && xPixel<265 && yPixel>=601 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=11 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=18 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=23 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=83 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=93 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=122 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=250 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=264 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=275 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=278 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=286 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=295 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=316 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=323 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=341 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=355 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=360 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=367 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=394 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=419 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=425 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=434 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=443 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=452 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=457 && yPixel<463) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=465 && yPixel<492) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=496 && yPixel<505) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=507 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=516 && yPixel<534) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=541 && yPixel<563) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=265 && xPixel<266 && yPixel>=564 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=4 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=21 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=28 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=86 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=126 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=210 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=288 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=293 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=306 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=316 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=325 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=333 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=358 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=361 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=366 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=370 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=382 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=391 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=401 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=426 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=442 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=447 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=452 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=457 && yPixel<486) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=487 && yPixel<492) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=496 && yPixel<504) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=504 && yPixel<506) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=506 && yPixel<510) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=510 && yPixel<518) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=519 && yPixel<524) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=524 && yPixel<527) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=534 && yPixel<542) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=542 && yPixel<562) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=563 && yPixel<571) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=266 && xPixel<267 && yPixel>=573 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=28 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=30 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=39 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=83 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=131 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=237 && yPixel<266) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=268 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=274 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=287 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=303 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b10000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=363 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=370 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=394 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=413 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=457 && yPixel<495) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=496 && yPixel<500) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=501 && yPixel<504) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=504 && yPixel<506) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=506 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=511 && yPixel<543) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=547 && yPixel<561) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=267 && xPixel<268 && yPixel>=574 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=1 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=3 && yPixel<5) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=7 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=34 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=35 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=37 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=42 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=46 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=81 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=131 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=134 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=192 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=199 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=243 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=270 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=279 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=288 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=298 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=349 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=359 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=368 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=390 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=403 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=450 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=453 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=458 && yPixel<462) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=463 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=490 && yPixel<499) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=499 && yPixel<507) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=507 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=513 && yPixel<549) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=554 && yPixel<557) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=557 && yPixel<565) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=565 && yPixel<574) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=268 && xPixel<269 && yPixel>=584 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=10 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=35 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=37 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=45 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=53 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=57 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=60 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=81 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=133 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=201 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=207 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=221 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=226 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=229 && yPixel<246) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=247 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=269 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=281 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=287 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=340 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=353 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=358 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=366 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=385 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=389 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=402 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=407 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=414 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=425 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=450 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=458 && yPixel<462) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=465 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=485 && yPixel<490) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=497 && yPixel<506) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=506 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=513 && yPixel<549) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=550 && yPixel<559) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=561 && yPixel<578) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=581 && yPixel<586) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=269 && xPixel<270 && yPixel>=586 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=8 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=10 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=29 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=38 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=41 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=44 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=73 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=75 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=78 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=105 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=108 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=123 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=126 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=128 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=134 && yPixel<142) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=146 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=150 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=154 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=157 && yPixel<161) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=171 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=180 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=201 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=217 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=231 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=238 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=245 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=258 && yPixel<266) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=267 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=278 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=283 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=302 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=339 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=350 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=351 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=356 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=363 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=396 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=415 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=457 && yPixel<462) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=463 && yPixel<478) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=483 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=487 && yPixel<493) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=494 && yPixel<507) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=507 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=513 && yPixel<559) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=565 && yPixel<579) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=580 && yPixel<587) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=270 && xPixel<271 && yPixel>=587 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=18 && yPixel<22) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=24 && yPixel<32) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=32 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=39 && yPixel<41) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=41 && yPixel<79) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=79 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=84 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=100 && yPixel<142) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=150 && yPixel<171) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=171 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=186 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=192 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=200 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=204 && yPixel<208) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=209 && yPixel<212) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=212 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=231 && yPixel<237) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=237 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=243 && yPixel<263) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=267 && yPixel<277) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=297 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=313 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=341 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=345 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=359 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=365 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=376 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=379 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=380 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=388 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=398 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=422 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=427 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=433 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=436 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=448 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=456 && yPixel<464) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=471 && yPixel<474) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=474 && yPixel<477) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=485 && yPixel<508) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=513 && yPixel<585) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=271 && xPixel<272 && yPixel>=588 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=0 && yPixel<271) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=271 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=330 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=331 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=333 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=341 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=371 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=379 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=383 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=390 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=393 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=414 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=419 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=424 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=437 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=441 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=456 && yPixel<467) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=467 && yPixel<476) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=477 && yPixel<512) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=514 && yPixel<588) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=272 && xPixel<273 && yPixel>=594 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=0 && yPixel<263) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=264 && yPixel<268) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=269 && yPixel<271) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=271 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=290 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=303 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=321 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=325 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=347 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=357 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=360 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=391 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11111111,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=419 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=439 && yPixel<454) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=454 && yPixel<457) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=457 && yPixel<468) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=468 && yPixel<476) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=477 && yPixel<512) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=513 && yPixel<588) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=273 && xPixel<274 && yPixel>=588 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=0 && yPixel<268) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=268 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=296 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=310 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=350 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=361 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=368 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=383 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=397 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=401 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=413 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=429 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=440 && yPixel<468) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=468 && yPixel<511) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=512 && yPixel<585) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=274 && xPixel<275 && yPixel>=589 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=0 && yPixel<268) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=268 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=311 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=329 && yPixel<363) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=370 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=381 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=388 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=395 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=412 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=426 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=440 && yPixel<460) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=462 && yPixel<466) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=469 && yPixel<511) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=512 && yPixel<588) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=275 && xPixel<276 && yPixel>=588 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=0 && yPixel<268) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=268 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=317 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=323 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=330 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=405 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=407 && yPixel<412) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=414 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=424 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=440 && yPixel<469) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=469 && yPixel<527) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=528 && yPixel<588) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=276 && xPixel<277 && yPixel>=595 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=0 && yPixel<181) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=181 && yPixel<184) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=184 && yPixel<268) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=268 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=330 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=391 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=397 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=404 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=413 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=440 && yPixel<467) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=467 && yPixel<588) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=277 && xPixel<278 && yPixel>=594 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=0 && yPixel<183) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=184 && yPixel<266) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=266 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=276 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=301 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=317 && yPixel<384) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=384 && yPixel<391) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=391 && yPixel<395) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=395 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=403 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=412 && yPixel<422) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=423 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=442 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=445 && yPixel<467) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=470 && yPixel<549) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=550 && yPixel<552) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=553 && yPixel<589) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=278 && xPixel<279 && yPixel>=589 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=0 && yPixel<216) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=216 && yPixel<222) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=223 && yPixel<233) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=236 && yPixel<246) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=247 && yPixel<256) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=261 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=266 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=272 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=277 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=302 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=320 && yPixel<325) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=325 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=331 && yPixel<353) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=355 && yPixel<365) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=366 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=386 && yPixel<391) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=391 && yPixel<395) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=395 && yPixel<399) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=399 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=407 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=412 && yPixel<437) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=438 && yPixel<442) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=442 && yPixel<467) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=469 && yPixel<470) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=470 && yPixel<489) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=491 && yPixel<551) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=554 && yPixel<587) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=279 && xPixel<280 && yPixel>=587 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=0 && yPixel<215) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=215 && yPixel<219) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=219 && yPixel<221) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=221 && yPixel<226) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=227 && yPixel<239) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=243 && yPixel<246) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=247 && yPixel<256) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=259 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=262 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=273 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=277 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=302 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=321 && yPixel<325) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=325 && yPixel<353) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=355 && yPixel<369) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=369 && yPixel<372) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=372 && yPixel<386) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=390 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=393 && yPixel<399) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=399 && yPixel<403) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=405 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=407 && yPixel<413) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=414 && yPixel<437) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=438 && yPixel<442) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=442 && yPixel<456) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=462 && yPixel<476) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=476 && yPixel<489) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=492 && yPixel<551) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=556 && yPixel<587) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=280 && xPixel<281 && yPixel>=587 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=0 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=64 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=67 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=95 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=108 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=109 && yPixel<220) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=222 && yPixel<226) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=227 && yPixel<232) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=233 && yPixel<244) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=245 && yPixel<260) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=262 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=276 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=279 && yPixel<285) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=287 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=306 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=311 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=332 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=338 && yPixel<351) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=351 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=359 && yPixel<403) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=404 && yPixel<413) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=417 && yPixel<432) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=436 && yPixel<440) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=440 && yPixel<455) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=464 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=512 && yPixel<538) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=539 && yPixel<553) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=553 && yPixel<558) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=561 && yPixel<566) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=568 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=602 && yPixel<612) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=612 && yPixel<622) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=281 && xPixel<282 && yPixel>=622 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=26 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=135 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=141 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=145 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=150 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=158 && yPixel<167) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=170 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=178 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=184 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=190 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=230 && yPixel<236) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=242 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=248 && yPixel<250) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=250 && yPixel<254) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=255 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=262 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=264 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=267 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=285 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=298 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=312 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=320 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=331 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=347 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=362 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=364 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=368 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=383 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=392 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=409 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=428 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=432 && yPixel<492) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=493 && yPixel<506) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=507 && yPixel<511) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=511 && yPixel<514) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=514 && yPixel<518) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=519 && yPixel<527) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=528 && yPixel<559) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=559 && yPixel<565) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=565 && yPixel<579) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=580 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=282 && xPixel<283 && yPixel>=608 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=2 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=3 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=25 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=28 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=31 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=167 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=229 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=241 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=265 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=323 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=328 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=333 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=343 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=428 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=431 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=440 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=442 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=453 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=457 && yPixel<463) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=466 && yPixel<537) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=541 && yPixel<551) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=554 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=569 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=283 && xPixel<284 && yPixel>=602 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=6 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=15 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=23 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=170 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=182 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=214 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=242 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=248 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=254 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=300 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=311 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=320 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=326 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=332 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=358 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=441 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=453 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=457 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=466 && yPixel<478) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=478 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=496 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=533 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=554 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=567 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=606 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=284 && xPixel<285 && yPixel>=615 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=2 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=3 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=6 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=14 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=16 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=20 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=23 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=32 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=164 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=168 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=217 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=240 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=253 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=262 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=323 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=330 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=350 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=360 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=433 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=460 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=473 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=477 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=483 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=485 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=491 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=498 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=500 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=504 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=513 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=518 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=525 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=529 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=536 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=541 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=567 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=576 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=590 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=600 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=605 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=610 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=285 && xPixel<286 && yPixel>=620 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=2 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=6 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=9 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=13 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=31 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=38 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=43 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=48 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=71 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=79 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=170 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=181 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=217 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=225 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=249 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=256 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=300 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=310 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=314 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=320 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=395 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=409 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=414 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=421 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=432 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=439 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=460 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=485 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=497 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=501 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=504 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=513 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=554 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=566 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=579 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=585 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=602 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=615 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=286 && xPixel<287 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=1 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=14 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=28 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=31 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=34 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=43 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=48 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=61 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=63 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=68 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=83 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=86 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=94 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=171 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=176 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=184 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=249 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=252 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=258 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=270 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=274 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=279 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=294 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=302 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=311 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=318 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=392 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=396 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=426 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=436 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=439 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=468 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=472 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=475 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=481 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=483 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=487 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=499 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=502 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=505 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=512 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=517 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=525 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=543 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=550 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=552 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=556 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=568 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=583 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=602 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=615 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=287 && xPixel<288 && yPixel>=625 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=6 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=8 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=13 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=34 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=38 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=82 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=85 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=88 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=96 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=154 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=180 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=183 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=186 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=188 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=202 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=205 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=215 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=245 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=271 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=289 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=301 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=309 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=318 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=388 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=417 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=427 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=434 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=438 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=457 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=468 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=474 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=481 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=483 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=489 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=506 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=515 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=517 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=523 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=537 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=543 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=582 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=603 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=624 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=288 && xPixel<289 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=7 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=15 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=20 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=25 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=28 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=32 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=38 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=66 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=69 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=76 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=78 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=83 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=86 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=91 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=100 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=103 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=108 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=110 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=157 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=165 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=170 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=178 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=190 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=199 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=210 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=215 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=228 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=237 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=243 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=253 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=269 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=302 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=304 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=318 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=376 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=386 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=398 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=402 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=412 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=423 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=426 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=433 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=441 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=462 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=466 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=468 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=472 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=475 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=482 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=494 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=515 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=519 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=522 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=528 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=540 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=549 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=561 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=575 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=584 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=608 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=289 && xPixel<290 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=7 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=25 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=31 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=34 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=41 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=46 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=50 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=53 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=60 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=69 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=71 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=82 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=98 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=102 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=106 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=107 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=176 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=183 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=187 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=199 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=202 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=217 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=224 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=239 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=246 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=248 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=252 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=256 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=261 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=266 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=268 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=277 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=301 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=312 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=317 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=383 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=385 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=393 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=404 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=409 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=418 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=427 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=431 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=436 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=453 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=457 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=468 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=472 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=476 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=478 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=490 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=495 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=498 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=500 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=516 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=522 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=529 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=533 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=541 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=558 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=568 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=574 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=587 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=609 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=625 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=290 && xPixel<291 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=4 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=7 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=16 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=28 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=37 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=75 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=77 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=79 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=81 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=174 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=182 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=193 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=207 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=215 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=219 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=231 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=237 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=242 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=261 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=266 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=280 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=295 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=315 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=327 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=334 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=394 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=397 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=411 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=419 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=426 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=435 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=450 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=457 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=469 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=474 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=476 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=478 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=488 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=498 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=505 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=511 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=524 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=528 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=532 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=534 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=542 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=558 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=562 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=567 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=598 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=606 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=627 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=291 && xPixel<292 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=5 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=7 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=12 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=20 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=34 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=82 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=154 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=156 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=169 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=182 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=184 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=187 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=193 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=198 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=212 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=217 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=221 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=224 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=244 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=248 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=251 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=268 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=276 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=283 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=302 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=307 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=317 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=324 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=330 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=340 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=347 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=376 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=379 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=383 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=384 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=394 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=398 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=405 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=418 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=430 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=442 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=447 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=455 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=463 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=475 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=479 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=484 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=492 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=496 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=513 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=525 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=530 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=532 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=540 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=551 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=557 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=563 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=577 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=588 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=608 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=292 && xPixel<293 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=2 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=25 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=29 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=33 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=71 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=104 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=170 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=176 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=182 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=188 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=215 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=225 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=241 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=246 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=254 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=265 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=274 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=295 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=298 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=303 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=314 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=319 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=327 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=386 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=390 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=393 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=398 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=414 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=418 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=437 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=450 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=457 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=463 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=469 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=472 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=477 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=485 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=496 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=503 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=524 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=530 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=543 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=551 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=568 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=583 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=598 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=609 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=293 && xPixel<294 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=0 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=23 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=32 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=35 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=41 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=44 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=52 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=55 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=59 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=63 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=72 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=74 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=78 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=81 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=93 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=101 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=105 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=169 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=175 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=181 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=185 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=192 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=198 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=214 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=224 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=231 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=233 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=242 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=255 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=257 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=262 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=271 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=274 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=285 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=300 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=312 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=391 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=393 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=398 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=411 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=433 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=438 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=457 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=460 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=462 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=471 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=475 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=494 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=499 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=503 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=508 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=521 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=526 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=545 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=550 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=571 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=584 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=595 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=618 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=294 && xPixel<295 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=2 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=3 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=6 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=10 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=18 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=21 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=27 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=30 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=35 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=39 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=51 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=76 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=83 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=92 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=155 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=158 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=173 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=180 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=190 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=196 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=204 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=212 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=219 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=226 && yPixel<235) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=243 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=249 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=253 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=256 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=262 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=266 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=268 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=272 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=292 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=300 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=308 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=316 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=328 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=389 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=391 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=394 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=403 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=413 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=422 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=427 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=441 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=462 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=465 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=471 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=476 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=482 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=494 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=499 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=503 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=511 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=517 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=524 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=534 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=539 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=546 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=552 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=556 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=571 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=586 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=592 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=600 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=604 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=611 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=623 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=295 && xPixel<296 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=4 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=8 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=21 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=28 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=31 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=76 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=79 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=152 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=154 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=176 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=181 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=186 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=249 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=252 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=263 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=280 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=289 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=310 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=313 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=321 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=337 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=344 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=351 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=392 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=416 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=423 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=440 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=443 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=448 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=455 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=459 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=469 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=490 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=503 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=505 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=519 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=527 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=531 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=543 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=559 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=580 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=597 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=610 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=614 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=296 && xPixel<297 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=4 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=11 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=19 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=26 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=82 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=87 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=91 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=168 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=219 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=231 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=243 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=250 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=255 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=259 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=265 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=277 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=288 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=295 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=300 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=310 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=321 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=332 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=347 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=406 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=412 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=420 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=433 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=448 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=451 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=453 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=461 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=473 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=481 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=495 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=511 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=523 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=530 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=542 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=544 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=559 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=578 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=586 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=597 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=605 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=611 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=297 && xPixel<298 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=6 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=13 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=17 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=22 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=40 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=82 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=90 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=100 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=104 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=107 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=109 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=163 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=172 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=176 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=184 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=197 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=216 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=241 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=245 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=248 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=257 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=264 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=283 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=285 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=293 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=302 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=306 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=317 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=323 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=347 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=356 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=371 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=374 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=386 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=398 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=420 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=427 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=436 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=459 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=463 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=472 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=477 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=479 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=484 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=496 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=498 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=500 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=502 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=505 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=508 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=513 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=537 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=542 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=564 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=580 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=592 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=605 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=614 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=624 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=632 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=298 && xPixel<299 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=24 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=28 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=36 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=68 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=78 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=79 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=89 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=97 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=113 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=116 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=170 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=178 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=184 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=209 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=217 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=242 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=249 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=252 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=258 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=261 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=274 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=293 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=305 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=318 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=333 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=338 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=348 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=413 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=426 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=439 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=442 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=469 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=474 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=480 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=483 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=485 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=494 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=502 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=504 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=528 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=534 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=541 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=554 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=566 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=580 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=585 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=590 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=594 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=604 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=614 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=626 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=299 && xPixel<300 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=0 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=33 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=51 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=56 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=63 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=70 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=83 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=90 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=95 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=116 && yPixel<117) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=117 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=160 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=172 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=179 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=187 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=193 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=195 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=208 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=218 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=239 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=250 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=255 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=259 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=268 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=270 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=279 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=293 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=298 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=311 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=317 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=325 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=334 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=340 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=347 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=354 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=378 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=394 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=399 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=409 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=417 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=423 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=429 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=440 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=447 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=449 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=451 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=454 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=458 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=461 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=470 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=482 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=497 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=514 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=519 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=529 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=531 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=535 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=545 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=568 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=577 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=589 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=591 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=594 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=608 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=300 && xPixel<301 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=18 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=34 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=47 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=64 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=69 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=73 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=82 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=87 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=92 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=98 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=100 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=170 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=175 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=180 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=210 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=216 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=235 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=246 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=255 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=264 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=267 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=276 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=284 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=298 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=303 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=312 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=317 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=324 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=336 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=347 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=349 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=370 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=371 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=398 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=414 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=418 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=421 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=424 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=433 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=435 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=455 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=459 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=467 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=473 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=483 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=490 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=497 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=506 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=521 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=538 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=545 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=554 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=580 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=613 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=630 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=301 && xPixel<302 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=12 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=18 && yPixel<21) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=23 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=31 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=67 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=73 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=75 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=78 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=164 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=179 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=186 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=191 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=201 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=209 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=213 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=244 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=247 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=256 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=273 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=299 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=305 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=310 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=319 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=324 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=331 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=342 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=349 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=412 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=417 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=434 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=441 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=448 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=462 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=471 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=473 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=477 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=483 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=485 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=497 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=513 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=515 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=524 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=531 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=538 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=545 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=550 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=568 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=577 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=585 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=604 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=611 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=616 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=302 && xPixel<303 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=0 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=45 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=75 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=90 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=98 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=101 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=105 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=110 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=157 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=173 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=176 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=194 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=230 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=237 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=249 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=253 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=259 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=263 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=268 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=270 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=275 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=293 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=300 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=321 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=339 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=410 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=418 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=435 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=442 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=447 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=450 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=460 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=471 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=474 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=486 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=492 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=505 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=514 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=530 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=535 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=538 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=554 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=561 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=568 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=591 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=599 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=609 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=614 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=619 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=629 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=303 && xPixel<304 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=21 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=28 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=33 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=75 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=80 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=149 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=162 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=185 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=188 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=194 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=201 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=206 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=217 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=241 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=246 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=255 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=257 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=272 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=276 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=291 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=309 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=315 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=323 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=330 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=339 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=375 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=409 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=417 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=421 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=422 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=432 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=435 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=438 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=452 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=460 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=466 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=468 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=478 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=482 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=487 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=491 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=497 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=502 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=505 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=523 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=538 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=549 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=578 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=588 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=304 && xPixel<305 && yPixel>=618 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=35 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=72 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=83 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=92 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=96 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=103 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=118 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=119 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=158 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=160 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=178 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=188 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=217 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=234 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=246 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=249 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=256 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=305 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=319 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=324 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=331 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=339 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=348 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=351 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=390 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=411 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=443 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=461 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=475 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=482 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=491 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=498 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=502 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=509 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=514 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=518 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=522 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=530 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=537 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=549 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=560 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=569 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=612 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=625 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=305 && xPixel<306 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=0 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=15 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=19 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=62 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=85 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=121 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=123 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=133 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=138 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=154 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=158 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=183 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=188 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=230 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=233 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=243 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=252 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=277 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=294 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=312 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=319 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=325 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=337 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=365 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=439 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=459 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=472 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=476 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=487 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=496 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=514 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=519 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=525 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=532 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=551 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=558 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=575 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=591 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=606 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=612 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=630 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=306 && xPixel<307 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=0 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=28 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=34 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=57 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=64 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=66 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=82 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=85 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=90 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=95 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=98 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=105 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=108 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=123 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=125 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=133 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=142 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=152 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=155 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=159 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=169 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=172 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=175 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=182 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=217 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=242 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=248 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=252 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=261 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=271 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=279 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=293 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=302 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=305 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=327 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=332 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=365 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=369 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=413 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=420 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=425 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=438 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=448 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=451 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=456 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=463 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=476 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=478 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=485 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=493 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=498 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=509 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=516 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=525 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=529 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=535 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=562 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=565 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=574 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=580 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=585 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=593 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=307 && xPixel<308 && yPixel>=599 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=26 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=48 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=55 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=63 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=68 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=75 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=84 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=86 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=91 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=106 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=108 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=109 && yPixel<112) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=112 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=121 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=124 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=165 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=211 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=237 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=243 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=245 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=254 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=264 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=271 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=274 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=279 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=325 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=335 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=340 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=351 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=412 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=426 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=436 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=459 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=468 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=480 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=487 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=493 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=503 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=507 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=512 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=520 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=526 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=543 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=554 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=563 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=568 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=573 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=581 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=591 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=594 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=308 && xPixel<309 && yPixel>=610 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=9 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=10 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=12 && yPixel<18) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=19 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=23 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=33 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=39 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=49 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=51 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=53 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=60 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=72 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=80 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=89 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=102 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=106 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=107 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=113 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=116 && yPixel<117) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=117 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=118 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=147 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=153 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=169 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=180 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=186 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=189 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=210 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=220 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=237 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=243 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=247 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=250 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=257 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=266 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=277 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=302 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=306 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=328 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=332 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=345 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=391 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=412 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=417 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=429 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=440 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=458 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=465 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=474 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=475 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=483 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=488 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=499 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=503 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=539 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=543 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=551 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=561 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=567 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=595 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=606 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=309 && xPixel<310 && yPixel>=617 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=0 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=17 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=52 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=55 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=69 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=74 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=81 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=92 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=98 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=100 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=106 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=115 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=130 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=135 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=142 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=175 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=179 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=193 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=202 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=215 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=221 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=237 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=246 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=252 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=262 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=298 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=306 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=319 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=322 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=341 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=349 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=359 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=414 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=419 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=441 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=447 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=451 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=453 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=459 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=468 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=469 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=472 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=483 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=489 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=494 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=503 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=510 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=539 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=542 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=551 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=561 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=574 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=606 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=619 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=310 && xPixel<311 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=22 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=27 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=40 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=58 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=64 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=74 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=84 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=86 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=100 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=108 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=110 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=156 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=161 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=170 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=174 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=182 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=192 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=199 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=204 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=219 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=232 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=244 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=259 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=278 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=294 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=319 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=325 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=332 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=337 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=352 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=359 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=363 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=369 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=400 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=420 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=423 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=435 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=439 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=451 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=466 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=470 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=487 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=491 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=496 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=501 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=504 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=509 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=514 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=542 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=548 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=558 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=563 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=570 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=584 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=593 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=601 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=616 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=624 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=311 && xPixel<312 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=19 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=24 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=34 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=93 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=96 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=104 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=113 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=125 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=156 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=172 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=177 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=218 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=243 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=249 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=255 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=278 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=291 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=292 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=320 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=348 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=359 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=439 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=455 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=469 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=475 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=481 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=483 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=497 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=501 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=547 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=551 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=559 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=570 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=583 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=588 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=604 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=611 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=614 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=626 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=312 && xPixel<313 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=0 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=24 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=29 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=34 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=37 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=41 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=45 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=50 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=61 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=70 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=95 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=109 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=118 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=145 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=152 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=158 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=168 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=171 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=194 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=209 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=215 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=229 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=237 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=241 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=243 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=251 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=255 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=270 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=295 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=300 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=326 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=348 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=361 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=366 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=402 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=414 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=426 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=429 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=441 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=449 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=463 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=469 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=473 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=481 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=495 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=506 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=510 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=514 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=524 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=574 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=593 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=615 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=313 && xPixel<314 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=0 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=44 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=50 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=57 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=64 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=67 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=69 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=89 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=92 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=99 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=105 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=110 && yPixel<119) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=119 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=122 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=124 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=150 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=154 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=157 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=175 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=177 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=191 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=202 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=205 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=219 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=230 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=237 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=244 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=249 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=251 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=269 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=275 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=290 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=300 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=302 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=304 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=305 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=327 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=333 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=346 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=363 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=403 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=409 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=417 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=432 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=435 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=446 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=452 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=458 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=473 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=482 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=491 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=506 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=513 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=531 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=537 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=541 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=551 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=562 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=570 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=589 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=610 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=619 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=314 && xPixel<315 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=34 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=38 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=45 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=47 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=52 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=67 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=78 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=85 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=88 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=105 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=114 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=132 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=144 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=149 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=153 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=158 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=170 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=191 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=193 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=197 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=201 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=209 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=225 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=235 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=244 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=252 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=254 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=263 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=274 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=302 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=327 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=340 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=362 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=368 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=370 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=374 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=383 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=390 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=416 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=420 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=431 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=440 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=444 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=464 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=472 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=481 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=491 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=499 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=513 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=517 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=524 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=528 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=535 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=542 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=552 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=556 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=569 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=572 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=589 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=597 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=611 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=623 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=629 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=315 && xPixel<316 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=9 && yPixel<19) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=19 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=24 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=28 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=33 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=49 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=61 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=68 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=75 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=77 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=108 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=111 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=112 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=144 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=150 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=174 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=192 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=208 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=212 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=216 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=234 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=245 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=253 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=267 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=336 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=341 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=353 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=359 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=376 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=388 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=392 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=405 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=408 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=425 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=429 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=440 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=445 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=463 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=469 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=472 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=476 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=486 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=492 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=494 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=518 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=525 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=531 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=535 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=559 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=562 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=603 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=609 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=618 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=316 && xPixel<317 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=12 && yPixel<25) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=31 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=43 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=45 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=50 && yPixel<86) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=87 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=90 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=101 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=108 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=158 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=176 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=186 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=190 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=200 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=210 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=223 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=236 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=246 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=251 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=253 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=261 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=295 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=303 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=354 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=361 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=382 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=394 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=405 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=408 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=418 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=431 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=441 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=452 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=459 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=476 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=481 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=493 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=503 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=514 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=530 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=538 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=585 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=595 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=618 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=317 && xPixel<318 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=30 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=33 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=37 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=42 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=50 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=52 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=69 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=72 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=75 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=104 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=106 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=107 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=111 && yPixel<112) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=112 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=117 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=118 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=122 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=126 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=127 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=130 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=137 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=144 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=155 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=173 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=193 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=196 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=219 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=223 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=226 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=231 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=250 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=255 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=258 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=264 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=287 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=291 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=296 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=301 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=315 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=337 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=346 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=355 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=364 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=394 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=415 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=420 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=428 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=442 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=454 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=463 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=469 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=477 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=487 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=512 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=526 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=530 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=537 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=549 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=579 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=584 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=592 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=611 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=614 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=620 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=318 && xPixel<319 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=34 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=39 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=51 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=62 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=65 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=69 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=110 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=111 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=114 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=119 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=124 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=144 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=149 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=150 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=156 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=162 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=172 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=177 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=193 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=199 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=209 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=212 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=233 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=243 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=267 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=276 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=299 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=321 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=334 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=340 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=342 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=344 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=346 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=371 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=377 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=386 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=404 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=409 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=422 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=426 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=443 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=450 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=473 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=476 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=480 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=491 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=493 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=498 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=501 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=504 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=512 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=521 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=560 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=569 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=591 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=597 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=623 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=629 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=319 && xPixel<320 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=24 && yPixel<26) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=26 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=31 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=40 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=51 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=60 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=72 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=85 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=90 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=100 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=106 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=121 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=124 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=126 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=139 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=159 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=164 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=177 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=195 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=203 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=208 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=219 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=230 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=240 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=244 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=248 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=254 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=255 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=263 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=265 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=271 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=277 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=297 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=319 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=322 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=333 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=334 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=343 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=352 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=358 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=391 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=398 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=404 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=413 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=420 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=423 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=431 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=441 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=446 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=448 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=462 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=474 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=529 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=553 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=562 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=571 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=585 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=605 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=619 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=622 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=320 && xPixel<321 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=32 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=37 && yPixel<39) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=41 && yPixel<44) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=44 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=52 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=55 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=68 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=72 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=85 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=87 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=100 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=107 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=111 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=119 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=123 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=142 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=162 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=167 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=177 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=188 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=214 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=225 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=236 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=246 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=253 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=285 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=300 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=318 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=348 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=373 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=375 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=383 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=405 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=415 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=432 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=435 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=437 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=442 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=445 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=459 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=467 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=472 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=481 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=490 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=495 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=513 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=520 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=530 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=544 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=553 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=571 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=579 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=603 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=611 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=321 && xPixel<322 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=0 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=17 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=24 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=34 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=36 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=41 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=52 && yPixel<65) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=66 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=71 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=74 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=76 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=84 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=91 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=106 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=110 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=115 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=121 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=127 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=133 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=135 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=145 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=169 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=171 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=177 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=182 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=190 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=193 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=200 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=209 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=220 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=238 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=246 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=248 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=254 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=257 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=258 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=263 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=266 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=274 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=287 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=289 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=293 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=298 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=301 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=319 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=329 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=370 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=393 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=403 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=411 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=415 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=430 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=435 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=446 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=461 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=466 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=472 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=478 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=488 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=512 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=515 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=522 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=526 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=535 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=540 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=545 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=550 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=553 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=558 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=572 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=581 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=593 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=598 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=322 && xPixel<323 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=18 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=21 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=35 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=38 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=43 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=53 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=71 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=89 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=116 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=122 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=127 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=132 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=143 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=148 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=171 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=178 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=191 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=209 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=218 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=238 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=245 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=249 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=254 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=269 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=276 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=282 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=289 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=299 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=312 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=333 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=346 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=363 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=369 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=377 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=381 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=384 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=396 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=407 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=417 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=433 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=435 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=445 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=466 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=472 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=506 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=510 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=512 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=520 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=529 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=536 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=546 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=550 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=553 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=562 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=575 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=584 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=596 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=323 && xPixel<324 && yPixel>=611 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=27 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=31 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=61 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=63 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=90 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=98 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=100 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=104 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=106 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=109 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=111 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=112 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=116 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=131 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=133 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=173 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=193 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=204 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=208 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=216 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=239 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=243 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=256 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=260 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=264 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=266 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=270 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=272 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=286 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=290 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=296 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=303 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=314 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=321 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=342 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=346 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=347 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=348 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=359 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=369 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=387 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=397 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=406 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=410 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=420 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=434 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=441 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=456 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=462 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=470 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=477 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=485 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=506 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=527 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=529 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=538 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=556 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=565 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=575 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=584 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=587 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=588 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=603 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=612 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=324 && xPixel<325 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=0 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=42 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=52 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=63 && yPixel<70) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=70 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=77 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=81 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=85 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=120 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=131 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=136 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=175 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=180 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=184 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=191 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=196 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=223 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=233 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=244 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=252 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=265 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=287 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=290 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=293 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=298 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=311 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=332 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=348 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=359 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=368 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=377 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=399 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=403 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=419 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=423 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=431 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=439 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=442 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=452 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=462 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=464 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=482 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=491 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=500 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=502 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=506 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=510 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=521 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=527 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=531 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=538 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=544 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=552 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=555 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=591 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=607 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=325 && xPixel<326 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=0 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=32 && yPixel<35) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=35 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=37 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=46 && yPixel<52) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=53 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=61 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=65 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=72 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=102 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=108 && yPixel<118) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=118 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=121 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=125 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=126 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=128 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=131 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=133 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=160 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=162 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=173 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=184 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=199 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=206 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=212 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=215 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=220 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=236 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=244 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=247 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=257 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=265 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=267 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=278 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=280 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=288 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=296 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=304 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=317 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=326 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=332 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=352 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=355 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=365 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=377 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=394 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=404 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=408 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=412 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=433 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=435 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=440 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=445 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=464 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=469 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=472 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=475 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=481 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=490 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=496 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=524 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=531 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=537 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=543 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=551 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=580 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=587 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=600 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=621 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=628 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=326 && xPixel<327 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=7 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=9 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=18 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=20 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=35 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=57 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=62 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=65 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=68 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=82 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=108 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=110 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=119 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=120 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=124 && yPixel<126) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=126 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=129 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=132 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=135 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=151 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=167 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=175 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=178 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=191 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=193 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=197 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=213 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=226 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=236 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=238 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=249 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=256 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=273 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=287 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=293 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=299 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=309 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=321 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=337 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=345 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=352 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=363 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=367 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=376 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=380 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=402 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=416 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=418 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=424 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=426 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=446 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=457 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=463 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=466 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=475 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=476 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=479 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=486 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=488 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=494 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=499 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=504 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=507 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=510 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=548 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=574 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=582 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=599 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=327 && xPixel<328 && yPixel>=613 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=0 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=33 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=59 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=65 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=67 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=69 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=85 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=105 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=107 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=122 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=131 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=138 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=147 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=182 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=189 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=195 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=203 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=214 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=230 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=236 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=239 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=248 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=267 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=275 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=286 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=301 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=338 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=345 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=356 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=364 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=380 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=404 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=406 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=411 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=418 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=423 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=433 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=443 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=448 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=455 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=463 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=464 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=468 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=474 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=486 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=491 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=495 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=498 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=504 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=509 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=525 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=531 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=548 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=560 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=574 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=594 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=600 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=614 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=328 && xPixel<329 && yPixel>=622 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=0 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=20 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=23 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=30 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=53 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=56 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=58 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=64 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=66 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=78 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=83 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=89 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=101 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=108 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=109 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=111 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=112 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=119 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=124 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=137 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=144 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=149 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=168 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=185 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=194 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=201 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=209 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=221 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=228 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=236 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=242 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=245 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=253 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=270 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=276 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=279 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=325 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=332 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=336 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=340 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=344 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=375 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=387 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=409 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=412 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=418 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=428 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=451 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=460 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=465 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=470 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=485 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=491 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=498 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=570 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=577 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=588 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=607 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=614 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=329 && xPixel<330 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=10 && yPixel<23) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=23 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=27 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=48 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=53 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=62 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=72 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=76 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=89 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=102 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=107 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=113 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=115 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=123 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=140 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=148 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=187 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=196 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=208 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=214 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=226 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=243 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=251 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=255 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=274 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=300 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=304 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=329 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=337 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=359 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=371 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=380 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=420 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=433 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=440 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=449 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=455 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=464 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=473 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=476 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=491 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=493 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=498 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=505 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=510 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=519 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=536 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=542 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=562 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=575 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=589 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=602 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=609 && yPixel<614) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=614 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=330 && xPixel<331 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=33 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=49 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=58 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=64 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=71 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=105 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=109 && yPixel<120) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=120 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=123 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=128 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=134 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=140 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=148 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=168 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=173 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=187 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=190 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=205 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=221 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=232 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=239 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=246 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=253 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=259 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=268 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=277 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=287 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=293 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=311 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=345 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=350 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=356 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=361 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=364 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=397 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=398 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=413 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=416 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=435 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=446 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=450 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=468 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=472 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=482 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=486 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=498 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=503 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=506 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=522 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=532 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=545 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=564 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=587 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=605 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=629 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=331 && xPixel<332 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=34 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=39 && yPixel<42) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=43 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=60 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=86 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=89 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=97 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=100 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=106 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=127 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=132 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=141 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=163 && yPixel<166) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=170 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=179 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=193 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=202 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=205 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=209 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=220 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=226 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=241 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=254 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=260 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=263 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=273 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=294 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=299 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=315 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=324 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=334 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=345 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=356 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=373 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=375 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=395 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=415 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=419 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=425 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=430 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=438 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=447 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=458 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=462 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=466 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=470 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=473 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=482 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=489 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=492 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=500 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=508 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=511 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=514 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=523 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=525 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=529 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=531 && yPixel<536) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=536 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=544 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=548 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=554 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=565 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=587 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=602 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=612 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=622 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=332 && xPixel<333 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=0 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=17 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=29 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=55 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=58 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=60 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=70 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=79 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=82 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=89 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=103 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=130 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=134 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=173 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=181 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=186 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=191 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=199 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=209 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=227 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=232 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=239 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=248 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=254 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=258 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=267 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=274 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=288 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=296 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=302 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=329 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=339 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=364 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=394 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=395 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=400 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=408 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=418 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=425 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=436 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=445 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=449 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=463 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=468 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=475 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=478 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=482 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=484 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=486 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=491 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=508 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=521 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=525 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=529 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=543 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=557 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=562 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=566 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=571 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=579 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=585 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=588 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=600 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=604 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=618 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=333 && xPixel<334 && yPixel>=623 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=0 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=29 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=54 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=56 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=60 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=79 && yPixel<82) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=83 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=105 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=108 && yPixel<123) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=123 && yPixel<125) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=125 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=128 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=131 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=181 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=188 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=198 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=202 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=204 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=216 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=226 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=231 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=237 && yPixel<241) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=241 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=253 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=257 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=261 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=274 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=281 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=299 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=311 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=314 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=320 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=341 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=360 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=363 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=370 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=375 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=378 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=382 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=387 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=394 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=407 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=414 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=415 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=420 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=428 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=443 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=453 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=461 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=474 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=482 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=490 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=497 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=500 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=506 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=508 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=513 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=523 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=526 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=545 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=560 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=564 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=574 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=577 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=589 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=608 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=618 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=334 && xPixel<335 && yPixel>=622 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=0 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=28 && yPixel<34) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=34 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=40 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=53 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=57 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=68 && yPixel<74) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=74 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=85 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=95 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=102 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=108 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=124 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=136 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=144 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=148 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=152 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=179 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=183 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=198 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=216 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=224 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=232 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=245 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=269 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=275 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=278 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=284 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=297 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=310 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=326 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=331 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=339 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=343 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=361 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=369 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=375 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=388 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=392 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=404 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=424 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=452 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=470 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=477 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=480 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=486 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=490 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=506 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=514 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=517 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=527 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=529 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=532 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=535 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=544 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=562 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=568 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=576 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=584 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=589 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=602 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=610 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=623 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=627 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=335 && xPixel<336 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=0 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=33 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=60 && yPixel<75) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=75 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=92 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=106 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=107 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=109 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=124 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=132 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=148 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=161 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=163 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=167 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=172 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=181 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=185 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=195 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=205 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=211 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=223 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=228 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=253 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=297 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=310 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=324 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=351 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=362 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=363 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=391 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=401 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=405 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=412 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=413 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=416 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=423 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=430 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=443 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=451 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=454 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=475 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=480 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=486 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=496 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=501 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=502 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=504 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=511 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=521 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=524 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=528 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=537 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=540 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=559 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=570 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=583 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=589 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=605 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=611 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=620 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=626 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=336 && xPixel<337 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=19 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=63 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=68 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=74 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=78 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=82 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=94 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=109 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=116 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=128 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=135 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=160 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=163 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=179 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=185 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=196 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=206 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=214 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=221 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=229 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=238 && yPixel<260) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=260 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=262 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=276 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=281 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=286 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=295 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=338 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=348 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=357 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=370 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=377 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=380 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=387 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=392 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=396 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=400 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=406 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=417 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=420 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=424 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=434 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=440 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=461 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=467 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=487 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=506 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=529 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=538 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=549 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=556 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=571 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=586 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=597 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=605 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=611 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=617 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=627 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=337 && xPixel<338 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=0 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=20 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=62 && yPixel<64) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=65 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=73 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=81 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=87 && yPixel<88) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=88 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=117 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=134 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=145 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=155 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=161 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=166 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=181 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=198 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=219 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=231 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=244 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=266 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=282 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=287 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=291 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=303 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=320 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=323 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=325 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=336 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=345 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=358 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=368 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=373 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=376 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=392 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=395 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=403 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=430 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=454 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=457 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=458 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=459 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=464 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=468 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=471 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=475 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=481 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=485 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=487 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=516 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=528 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=538 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=542 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=571 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=586 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=590 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=600 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=606 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=627 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=338 && xPixel<339 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=0 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=23 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=54 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=58 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=70 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=80 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=97 && yPixel<100) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=101 && yPixel<120) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=120 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=126 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=127 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=128 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=134 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=139 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=146 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=158 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=175 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=183 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=185 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=191 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=194 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=204 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=215 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=230 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=233 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=243 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=251 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=258 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=276 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=290 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=308 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=315 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=320 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=325 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=327 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=338 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=347 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=352 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=368 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=375 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=379 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=386 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=392 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=398 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=406 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=422 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=425 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=450 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=465 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=467 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=481 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=492 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=495 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=517 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=526 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=533 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=537 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=552 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=557 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=568 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=578 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=586 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=598 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=607 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=620 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=625 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=339 && xPixel<340 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=0 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=25 && yPixel<38) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=38 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=45 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=63 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=77 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=80 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=97 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=101 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=106 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=109 && yPixel<121) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=121 && yPixel<128) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=131 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=149 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=186 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=193 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=197 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=202 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=208 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=217 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=230 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=250 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=259 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=263 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=271 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=277 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=285 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=288 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=290 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=301 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=308 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=318 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=325 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=328 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=336 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=352 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=369 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=371 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=374 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=381 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=397 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=409 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=417 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=452 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=458 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=461 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=465 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=478 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=488 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=495 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=496 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=513 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=525 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=527 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=533 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=543 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=552 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=569 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=575 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=582 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=606 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=612 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=629 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=340 && xPixel<341 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=22 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=37 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=52 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=61 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=72 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=76 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=80 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=82 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=85 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=94 && yPixel<97) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=100 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=107 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=126 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=141 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=147 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=188 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=192 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=198 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=209 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=227 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=232 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=238 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=252 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=256 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=262 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=269 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=286 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=295 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=307 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=315 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=320 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=323 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=327 && yPixel<333) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=333 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=335 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=345 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=358 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=367 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=373 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=376 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=390 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=395 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=401 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=409 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=419 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=421 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=436 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=443 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=451 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=463 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=465 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=478 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=483 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=484 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=498 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=513 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=525 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=534 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=537 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=545 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=558 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=562 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=576 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=581 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=593 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=604 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=619 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=341 && xPixel<342 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=14 && yPixel<29) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=31 && yPixel<41) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=41 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=57 && yPixel<72) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=72 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=76 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=95 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=103 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=118 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=132 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=166 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=169 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=173 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=178 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=187 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=192 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=198 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=209 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=213 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=219 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=227 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=232 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=237 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=248 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=251 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=257 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=261 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=269 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=276 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=291 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=297 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=303 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=308 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=320 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=333 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=341 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=347 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=357 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=362 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=366 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=373 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=383 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=391 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=404 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=412 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=418 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=426 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=437 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=451 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=458 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=467 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=474 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=498 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=536 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=537 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=550 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=556 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=559 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=565 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=569 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=580 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=602 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=342 && xPixel<343 && yPixel>=614 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=19 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=32 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=38 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=42 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=44 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=58 && yPixel<71) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=71 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=81 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=101 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=107 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=119 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=131 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=156 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=170 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=180 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=184 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=186 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=201 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=207 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=219 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=225 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=231 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=244 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=267 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=276 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=286 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=300 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=322 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=323 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=328 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=336 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=348 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=358 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=367 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=373 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=391 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=395 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=402 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=412 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=415 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=417 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=426 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=428 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=434 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=443 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=450 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=461 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=470 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=474 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=481 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=488 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=497 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=508 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=514 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=539 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=547 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=555 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=574 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=587 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=595 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=613 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=621 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=343 && xPixel<344 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=22 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=36 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=46 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=48 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=55 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=67 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=71 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=78 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=92 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=98 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=105 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=107 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=112 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=121 && yPixel<127) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=127 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=137 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=140 && yPixel<142) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=142 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=153 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=156 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=162 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=176 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=187 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=196 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=209 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=224 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=229 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=232 && yPixel<247) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=248 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=254 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=268 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=277 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=286 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=304 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=317 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=331 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=336 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=347 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=359 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=386 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=392 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=395 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=409 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=418 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=443 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=450 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=452 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=459 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=471 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=474 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=481 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=499 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=504 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=507 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=525 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=556 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=557 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=563 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=572 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=582 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=592 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=600 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=615 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=344 && xPixel<345 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=14 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=17 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=21 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=45 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=50 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=63 && yPixel<80) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=80 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=94 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=101 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=105 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=106 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=109 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=115 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=117 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=158 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=170 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=180 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=199 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=231 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=243 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=250 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=255 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=268 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=272 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=277 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=286 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=296 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=298 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=302 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=310 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=316 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=320 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=329 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=335 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=339 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=366 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=370 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=372 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=379 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=384 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=395 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=399 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=414 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=430 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=440 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=449 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=458 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=460 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=461 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=464 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=465 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=466 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=475 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=478 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=481 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=486 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=501 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=509 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=519 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=524 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=530 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=533 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=534 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=537 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=553 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=558 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=565 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=580 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=589 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=602 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=618 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=628 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=345 && xPixel<346 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=11 && yPixel<17) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=17 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=22 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=49 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=62 && yPixel<71) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=72 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=79 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=90 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=103 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=105 && yPixel<107) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=107 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=112 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=128 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=131 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=145 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=149 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=172 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=177 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=186 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=216 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=222 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=231 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=233 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=236 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=246 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=267 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=271 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=278 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=294 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=298 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=302 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=307 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=324 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=330 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=333 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=349 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=360 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=366 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=371 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=403 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=417 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=432 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=440 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=452 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=460 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=467 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=480 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=482 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=491 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=494 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=496 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=504 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=532 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=550 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=571 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=580 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=589 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=598 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=346 && xPixel<347 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=0 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=25 && yPixel<32) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=32 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=39 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=61 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=66 && yPixel<72) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=72 && yPixel<74) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=74 && yPixel<79) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=79 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=94 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=104 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=108 && yPixel<120) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=120 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=138 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=144 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=150 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=179 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=182 && yPixel<184) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=184 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=190 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=204 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=221 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=225 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=238 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=247 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=257 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=262 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=279 && yPixel<282) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=282 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=284 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=289 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=303 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=307 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=313 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=331 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=336 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=341 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=357 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=368 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=384 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=390 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=395 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=400 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=409 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=417 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=422 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=430 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=446 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=453 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=461 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=467 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=469 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=478 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=481 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=499 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=503 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=506 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=509 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=510 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=512 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=513 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=514 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=536 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=549 && yPixel<555) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=555 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=562 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=577 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=584 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=597 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=617 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=347 && xPixel<348 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=0 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=28 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=53 && yPixel<66) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=66 && yPixel<77) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=77 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=80 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=86 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=91 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=112 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=126 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=135 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=146 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=176 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=182 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=189 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=196 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=205 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=232 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=247 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=264 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=272 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=280 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=296 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=302 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=318 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=322 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=325 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=336 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=356 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=359 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=363 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=368 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=377 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=380 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=392 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=400 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=403 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=406 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=410 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=426 && yPixel<435) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=435 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=438 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=452 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=474 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=477 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=485 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=491 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=493 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=500 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=504 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=515 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=517 && yPixel<523) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=523 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=528 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=536 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=541 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=551 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=559 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=562 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=571 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=580 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=586 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=603 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=608 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=612 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=625 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=348 && xPixel<349 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=0 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=28 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=51 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=58 && yPixel<68) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=68 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=97 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=102 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=104 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=109 && yPixel<111) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=111 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=129 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=132 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=137 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=144 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=149 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=153 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=177 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=189 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=193 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=199 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=207 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=219 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=222 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=237 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=252 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=285 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=294 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=304 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=344 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=349 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=354 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=359 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=365 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=369 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=371 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=380 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=382 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=410 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=414 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=420 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=434 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=443 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=447 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=452 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=466 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=476 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=492 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=497 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=504 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=506 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=510 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=513 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=517 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=536 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=541 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=549 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=553 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=556 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=565 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=584 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=593 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=609 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=623 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=349 && xPixel<350 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=0 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=28 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=49 && yPixel<53) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=53 && yPixel<58) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=58 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=63 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=78 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=95 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=110 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=140 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=150 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=155 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=184 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=194 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=198 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=201 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=206 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=219 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=225 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=237 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=268 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=272 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=300 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=315 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=322 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=344 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=359 && yPixel<364) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=364 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=368 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=386 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=412 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=419 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=430 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=443 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=449 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=462 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=465 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=475 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=497 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=503 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=508 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=519 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=528 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=532 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=539 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=540 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=546 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=552 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=555 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=557 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=570 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=604 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=609 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=624 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=630 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=350 && xPixel<351 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=0 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=30 && yPixel<48) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=48 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=54 && yPixel<57) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=58 && yPixel<76) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=76 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=80 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=99 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=105 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=119 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=156 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=168 && yPixel<172) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=172 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=175 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=184 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=185 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=198 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=204 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=222 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=231 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=240 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=247 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=269 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=289 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=314 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=321 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=325 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=335 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=341 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=347 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=358 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=371 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=378 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=388 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=397 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=410 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=446 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=452 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=458 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=466 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=491 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=515 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=519 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=522 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=533 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=546 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=557 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=571 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=602 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=351 && xPixel<352 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=2 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=13 && yPixel<16) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=16 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=36 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=47 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=57 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=60 && yPixel<63) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=63 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=67 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=94 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=102 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=109 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=112 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=156 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=169 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=200 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=208 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=223 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=241 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=249 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=266 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=270 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=292 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=299 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=304 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=309 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=329 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=342 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=373 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=384 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=388 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=399 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=402 && yPixel<409) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=409 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=418 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=429 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=435 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=443 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=450 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=471 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=483 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=488 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=493 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=501 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=520 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=552 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=568 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=573 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=586 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=590 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=594 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=600 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=603 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=613 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=352 && xPixel<353 && yPixel>=625 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=21 && yPixel<30) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=30 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=41 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=51 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=60 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=64 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=84 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=106 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=154 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=160 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=162 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=168 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=182 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=194 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=211 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=223 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=238 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=242 && yPixel<246) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=247 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=251 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=262 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=265 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=269 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=277 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=292 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=310 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=322 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=341 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=356 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=364 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=375 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=388 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=425 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=433 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=442 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=445 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=455 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=489 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=491 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=494 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=498 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=505 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=518 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=522 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=530 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=537 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=542 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=547 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=575 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=589 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=601 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=617 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=629 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=353 && xPixel<354 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=26 && yPixel<37) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=37 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=47 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=55 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=75 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=84 && yPixel<93) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=93 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=95 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=99 && yPixel<102) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=103 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=109 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=136 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=140 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=149 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=160 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=175 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=187 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=190 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=198 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=217 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=239 && yPixel<242) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=242 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=251 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=257 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=264 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=269 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=278 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=296 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=311 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=317 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=341 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=344 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=347 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=353 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=367 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=369 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=379 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=383 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=389 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=403 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=405 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=408 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=428 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=432 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=443 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=458 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=464 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=466 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=468 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=476 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=481 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=487 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=494 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=521 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=526 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=535 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=546 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=552 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b10000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=578 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=586 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=601 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=608 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=627 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=354 && xPixel<355 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=0 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=44 && yPixel<55) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=55 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=87 && yPixel<90) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=90 && yPixel<92) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=92 && yPixel<100) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=100 && yPixel<106) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=108 && yPixel<109) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=109 && yPixel<116) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=116 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=140 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=173 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=201 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=207 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=219 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=229 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=233 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=243 && yPixel<250) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=250 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=263 && yPixel<266) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=267 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=269 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=274 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=292 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=303 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=309 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=329 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=341 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=345 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=350 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=358 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=379 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=395 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=405 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=420 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=425 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=431 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=437 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=439 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=443 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=456 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=460 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=467 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=471 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=479 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=488 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=496 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=497 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=510 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=515 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=526 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=540 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=544 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=561 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=568 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=587 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=590 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=602 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=606 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=609 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=617 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=355 && xPixel<356 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=2 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=5 && yPixel<16) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=18 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=41 && yPixel<55) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=55 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=60 && yPixel<65) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=65 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=72 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=89 && yPixel<92) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=95 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=114 && yPixel<119) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=119 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=145 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=156 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=164 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=181 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=185 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=190 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=197 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=201 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=210 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=225 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=232 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=235 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=242 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=254 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=266 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=270 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=279 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=283 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=287 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=294 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=299 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=310 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=314 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=320 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=332 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=338 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=346 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=361 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=376 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=394 && yPixel<404) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=404 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=410 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=413 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=422 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=430 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=444 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=451 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=467 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=489 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=493 && yPixel<495) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=495 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=507 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=513 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=515 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=518 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=519 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=523 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=541 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=554 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=557 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=560 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=561 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=566 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=574 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=582 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=585 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=599 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=606 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=622 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=356 && xPixel<357 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=1 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=8 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=18 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=24 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=42 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=51 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=56 && yPixel<65) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=65 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=72 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=79 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=83 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=96 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=118 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=149 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=158 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=162 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=196 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=207 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=211 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=217 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=226 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=231 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=234 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=243 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=247 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=251 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=263 && yPixel<271) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=271 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=279 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=288 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=299 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=315 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=321 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=326 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=340 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=348 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=355 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=363 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=372 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=376 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=378 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=379 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=386 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=400 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=411 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=417 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=437 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=449 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=480 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=487 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=489 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=499 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=502 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=513 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=521 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=523 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=553 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=563 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=587 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=606 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=357 && xPixel<358 && yPixel>=628 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=4 && yPixel<16) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=16 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=19 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=40 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=44 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=49 && yPixel<67) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=67 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=73 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=83 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=89 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=103 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=152 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=158 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=163 && yPixel<167) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=167 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=170 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=182 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=183 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=192 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=204 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=214 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=221 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=226 && yPixel<246) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=246 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=248 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=255 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=261 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=280 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=291 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=315 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=335 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=344 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=351 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=357 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=359 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=371 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=392 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=393 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=396 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=412 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=422 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=424 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=433 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=438 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=443 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=483 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=494 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=519 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=522 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=529 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=554 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=562 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=576 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=583 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=598 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=606 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=609 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=617 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=358 && xPixel<359 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=0 && yPixel<22) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=22 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=25 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=38 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=41 && yPixel<67) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=68 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=71 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=96 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=105 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=154 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=160 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=169 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=180 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=181 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=191 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=197 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=204 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=212 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=215 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=222 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=228 && yPixel<244) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=245 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=257 && yPixel<265) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=265 && yPixel<275) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=275 && yPixel<281) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=281 && yPixel<289) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=289 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=297 && yPixel<300) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=302 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=311 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=323 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=326 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=331 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=339 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=348 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=363 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=368 && yPixel<373) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=373 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=389 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=396 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=399 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=401 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=406 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=418 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=421 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=426 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=433 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=437 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=499 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=501 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=509 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=512 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=514 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=515 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=517 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=518 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=523 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=531 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=534 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=550 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=562 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=572 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=589 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=596 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=604 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=615 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=621 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=359 && xPixel<360 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=0 && yPixel<25) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=25 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=40 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=44 && yPixel<64) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=65 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=68 && yPixel<91) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=98 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=102 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=107 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=137 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=155 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=165 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=186 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=192 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=197 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=203 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=217 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=221 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=240 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=244 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=248 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=250 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=252 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=259 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=277 && yPixel<280) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=280 && yPixel<283) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=283 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=289 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=300 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=309 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=315 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=330 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=343 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=349 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=356 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=360 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=362 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=371 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=393 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=397 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=405 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=419 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=434 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=445 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=455 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=457 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=461 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=467 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=481 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=498 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=509 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=514 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=517 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=535 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=553 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=571 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=579 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=604 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=622 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=626 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=360 && xPixel<361 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=28 && yPixel<30) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=30 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=39 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=41 && yPixel<47) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=49 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=56 && yPixel<62) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=63 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=65 && yPixel<68) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=68 && yPixel<71) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=71 && yPixel<89) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=89 && yPixel<92) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=94 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=103 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=107 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=110 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=148 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=153 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=166 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=188 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=196 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=205 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=208 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=223 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=249 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=252 && yPixel<263) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=263 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=273 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=278 && yPixel<281) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=281 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=287 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=289 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=318 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=339 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=358 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=373 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=379 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=392 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=425 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=435 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=446 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=451 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=464 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=487 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=497 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=512 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=524 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=531 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=542 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=547 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=558 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=561 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=575 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=585 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=589 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=593 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=600 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=611 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=616 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=361 && xPixel<362 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=6 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=20 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=22 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=24 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=35 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=50 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=55 && yPixel<64) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=64 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=73 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=81 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=90 && yPixel<102) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=102 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=135 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=140 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=149 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=165 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=191 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=196 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=202 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=219 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=224 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=238 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=247 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=251 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=270 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=277 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=281 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=291 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=294 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=297 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=313 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=320 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=324 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=328 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=334 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=340 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=354 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=355 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=361 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=367 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=390 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=392 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=406 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=422 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=431 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=445 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=452 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=463 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=471 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=476 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=491 && yPixel<492) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=492 && yPixel<501) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=501 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=505 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=508 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=515 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=523 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=529 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=535 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=538 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=560 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=568 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=609 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=362 && xPixel<363 && yPixel>=625 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=8 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=10 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=13 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=20 && yPixel<23) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=23 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=37 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=56 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=61 && yPixel<69) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=69 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=74 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=76 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=82 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=90 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=96 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=100 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=104 && yPixel<112) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=112 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=114 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=133 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=137 && yPixel<142) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=146 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=155 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=171 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=191 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=193 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=202 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=213 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=223 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=239 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=251 && yPixel<259) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=261 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=267 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=273 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=276 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=281 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=287 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=322 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=333 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=337 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=344 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=370 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=433 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=444 && yPixel<461) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=461 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=469 && yPixel<478) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=478 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=480 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=489 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=496 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=500 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=504 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=511 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=513 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=528 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=536 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=539 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=554 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=567 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=573 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=584 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=595 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=604 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=606 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=610 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=614 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=625 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=363 && xPixel<364 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=0 && yPixel<20) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=22 && yPixel<24) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=24 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=27 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=38 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=54 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=60 && yPixel<67) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=67 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=72 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=76 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=82 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=86 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=89 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=97 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=124 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=128 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=134 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=136 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=140 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=147 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=151 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=161 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=164 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=168 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=172 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=175 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=204 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=217 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=225 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=234 && yPixel<246) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=247 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=251 && yPixel<270) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=270 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=278 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=295 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=306 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=312 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=317 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=318 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=320 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=322 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=361 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=387 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=421 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=433 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=444 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=491 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=493 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=499 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=508 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=519 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=531 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=544 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=549 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=552 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=555 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=559 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=570 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=575 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=592 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=596 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=615 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=623 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=628 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=364 && xPixel<365 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=7 && yPixel<10) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=10 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=15 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=17 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=19 && yPixel<24) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=28 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=31 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=44 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=50 && yPixel<56) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=56 && yPixel<61) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=61 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=63 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=65 && yPixel<69) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=69 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=75 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=95 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=105 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=135 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=139 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=148 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=153 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=160 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=167 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=172 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=209 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=242 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=249 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=286 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=296 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=317 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=362 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=368 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=371 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=377 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=383 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=392 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=400 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=409 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=423 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=426 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=435 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=440 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=444 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=451 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=455 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=464 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=474 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=482 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=496 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=504 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=509 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=516 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=517 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=528 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=532 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=542 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=544 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=550 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=559 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=574 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=578 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=580 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=584 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=597 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=603 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=614 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=617 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=365 && xPixel<366 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=0 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=48 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=51 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=55 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=62 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=65 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=67 && yPixel<74) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=74 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=83 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=94 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=98 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=101 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=141 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=154 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=161 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=163 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=171 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=200 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=206 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=221 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=236 && yPixel<264) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=264 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=268 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=279 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=282 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=292 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=299 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=305 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=312 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=316 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=317 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=339 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=340 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=352 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=362 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=378 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=387 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=401 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=410 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=423 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=430 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=436 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=438 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=444 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=449 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=452 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=466 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=469 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=478 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=489 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=493 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=497 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=515 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=520 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=541 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=542 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=554 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=557 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=573 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=580 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=589 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=603 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=628 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=366 && xPixel<367 && yPixel>=630 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=5 && yPixel<20) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=20 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=48 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=66 && yPixel<71) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=78 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=101 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=149 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=162 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=176 && yPixel<180) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=180 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=190 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=197 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=201 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=207 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=213 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=231 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=233 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=243 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=251 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=263 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=281 && yPixel<286) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=286 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=287 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=300 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=311 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=314 && yPixel<317) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=319 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=330 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=345 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=352 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=357 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=380 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=383 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=387 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=399 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=410 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=416 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=421 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=425 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=428 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=432 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=437 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=442 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=444 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=448 && yPixel<451) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=452 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=460 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=470 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=480 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=481 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=482 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=486 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=488 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=489 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=493 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=505 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=509 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=514 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=521 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=534 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=538 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=549 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=564 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=582 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=607 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=613 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=633 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=367 && xPixel<368 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=9 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=49 && yPixel<55) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=56 && yPixel<71) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=71 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=77 && yPixel<79) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=79 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=99 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=105 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=118 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=148 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=154 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=165 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=183 && yPixel<185) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=185 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=187 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=220 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=226 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=231 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=233 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=243 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=283 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=288 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=301 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=313 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=320 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=324 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=325 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=327 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=330 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=338 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=355 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=358 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=362 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=372 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=380 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=389 && yPixel<395) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=395 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=407 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=409 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=420 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=430 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=433 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=444 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=455 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=458 && yPixel<479) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=479 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=482 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=487 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=488 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=491 && yPixel<510) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=510 && yPixel<515) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=515 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=526 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=530 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=534 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=540 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=548 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=552 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=560 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=576 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=580 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=596 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=601 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=606 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=623 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=635 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=368 && xPixel<369 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=0 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=40 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=55 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=65 && yPixel<71) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=71 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=97 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=108 && yPixel<113) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=113 && yPixel<118) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=118 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=148 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=157 && yPixel<161) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=163 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=180 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=183 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=187 && yPixel<189) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=194 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=206 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=214 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=239 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=249 && yPixel<253) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=253 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=288 && yPixel<297) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=297 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=301 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=310 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=311 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=315 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=326 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=339 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=349 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=364 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=373 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=374 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=379 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=385 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=388 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=392 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=407 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=432 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=436 && yPixel<442) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=446 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=449 && yPixel<455) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=455 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=462 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=481 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=486 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=493 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=502 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=508 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=514 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=523 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=534 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=540 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=548 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=555 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=576 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=579 && yPixel<591) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=596 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=614 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=618 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=622 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=369 && xPixel<370 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=6 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=39 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=42 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=48 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=58 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=67 && yPixel<69) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=69 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=72 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=77 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=94 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=108 && yPixel<111) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=111 && yPixel<112) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=112 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=117 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=137 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=142 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=147 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=153 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=163 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=176 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=179 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=183 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=187 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=190 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=204 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=218 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=227 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=229 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=233 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=238 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=243 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=247 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=250 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=253 && yPixel<261) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=262 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=269 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=293 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=305 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=307 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=310 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=317 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=319 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=323 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=335 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=342 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=352 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=353 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=361 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=365 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=377 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=401 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=411 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=416 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=421 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=433 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=443 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=455 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=459 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=480 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=524 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=534 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=554 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=562 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=576 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=582 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=587 && yPixel<591) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=597 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=607 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=613 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=615 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=618 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=625 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=627 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=370 && xPixel<371 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=0 && yPixel<20) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=20 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=26 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=47 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=51 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=55 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=57 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=61 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=70 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=75 && yPixel<84) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=84 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=92 && yPixel<97) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=97 && yPixel<101) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=102 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=110 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=136 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=147 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=154 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=157 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=160 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=165 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=206 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=218 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=226 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=237 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=256 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=276 && yPixel<289) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=289 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=291 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=303 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=307 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=310 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=320 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=328 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=335 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=358 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=363 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=367 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=386 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=389 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=395 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=409 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=419 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=443 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=447 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=456 && yPixel<458) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=458 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=481 && yPixel<493) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=493 && yPixel<496) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=496 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=525 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=528 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=535 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=541 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=548 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=565 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=572 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=588 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=599 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=604 && yPixel<609) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=611 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=615 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=371 && xPixel<372 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=0 && yPixel<13) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=13 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=25 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=29 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=30 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=32 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=43 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=47 && yPixel<58) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=58 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=62 && yPixel<67) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=67 && yPixel<78) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=78 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=93 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=98 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=106 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=107 && yPixel<109) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=109 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=150 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=154 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=156 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=166 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=170 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=178 && yPixel<189) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=189 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=201 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=208 && yPixel<223) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=223 && yPixel<242) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=242 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=270 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=275 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=277 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=282 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=304 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=308 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=310 && yPixel<313) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=313 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=323 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=328 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=339 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=356 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=372 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=374 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=380 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=389 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=393 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=410 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=412 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=437 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=441 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=443 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=472 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=478 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=517 && yPixel<528) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=528 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=534 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=540 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=547 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=570 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=590 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=594 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=603 && yPixel<605) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=605 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=612 && yPixel<613) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=613 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=614 && yPixel<619) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=623 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=372 && xPixel<373 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=0 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=39 && yPixel<49) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=50 && yPixel<57) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=57 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=88 && yPixel<95) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=96 && yPixel<99) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=99 && yPixel<102) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=102 && yPixel<103) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=103 && yPixel<107) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=107 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=150 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=165 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=187 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=198 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=201 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=215 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=227 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=238 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=264 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=269 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=280 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=287 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=291 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=294 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=303 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=311 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=318 && yPixel<323) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=323 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=332 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=335 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=344 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=349 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=374 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=376 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=383 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=387 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=403 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=431 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=443 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=449 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=456 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=461 && yPixel<469) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=469 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=480 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=504 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=514 && yPixel<537) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=537 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=543 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=544 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=555 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=572 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=582 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=593 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=609 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=612 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=616 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=624 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=373 && xPixel<374 && yPixel>=627 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=5 && yPixel<11) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=11 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=32 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=48 && yPixel<64) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=64 && yPixel<69) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=69 && yPixel<73) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=73 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=87 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=104 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=108 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=114 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=140 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=146 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=165 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=206 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=213 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=230 && yPixel<233) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=233 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=240 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=248 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=268 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=275 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=277 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=281 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=285 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=293 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=298 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=302 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=309 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=332 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=339 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=345 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=353 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=356 && yPixel<365) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=365 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=377 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=387 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=391 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=406 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=412 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=432 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=438 && yPixel<441) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=443 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=446 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=457 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=469 && yPixel<474) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=474 && yPixel<488) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=488 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=504 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=512 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=532 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=536 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=555 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=567 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=569 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=595 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=619 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=374 && xPixel<375 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=5 && yPixel<7) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=7 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=18 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=20 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=32 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=40 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=64 && yPixel<70) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=70 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=74 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=99 && yPixel<104) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=105 && yPixel<108) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=108 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=110 && yPixel<115) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=115 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=147 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=152 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=166 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=195 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=204 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=206 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=221 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=226 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=232 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=270 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=284 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=292 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=297 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=302 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=318 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=329 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=332 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=338 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=340 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=341 && yPixel<346) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=346 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=350 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=357 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=362 && yPixel<370) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=370 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=378 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=384 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=389 && yPixel<398) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=398 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=402 && yPixel<406) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=406 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=414 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=439 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=445 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=470 && yPixel<484) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=484 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=485 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=494 && yPixel<497) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=497 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=506 && yPixel<512) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=512 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=524 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=532 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=543 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=547 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=549 && yPixel<557) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=557 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=559 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=565 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=579 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=588 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=590 && yPixel<591) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=591 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=599 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=612 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=625 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=375 && xPixel<376 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=8 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=14 && yPixel<15) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=15 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=17 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=20 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=22 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=51 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=68 && yPixel<78) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=78 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=97 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=103 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=107 && yPixel<110) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=110 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=146 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=164 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=211 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=218 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=232 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=238 && yPixel<252) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=252 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=261 && yPixel<264) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=265 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=270 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=277 && yPixel<289) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=289 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=294 && yPixel<298) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=303 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=305 && yPixel<306) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=306 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=312 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=323 && yPixel<325) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=325 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=334 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=341 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=344 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=349 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=356 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=384 && yPixel<389) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=389 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=390 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=404 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=409 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=425 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=445 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=498 && yPixel<502) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=502 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=503 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=505 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=513 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=524 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=530 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=558 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=592 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=602 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=608 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=611 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=617 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=376 && xPixel<377 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=14 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=17 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=19 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=27 && yPixel<36) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=36 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=46 && yPixel<50) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=51 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=53 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=55 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=62 && yPixel<78) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=78 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=105 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=128 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=134 && yPixel<143) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=143 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=146 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=155 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=156 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=164 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=213 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=225 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=229 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=236 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=258 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=259 && yPixel<263) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=263 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=276 && yPixel<297) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=297 && yPixel<301) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=301 && yPixel<302) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=302 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=306 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=309 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=316 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=321 && yPixel<325) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=325 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=334 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=335 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=346 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=348 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=352 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=378 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=409 && yPixel<426) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=426 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=439 && yPixel<443) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=453 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=454 && yPixel<466) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=466 && yPixel<479) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=479 && yPixel<480) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=480 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=504 && yPixel<507) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=507 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=508 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=509 && yPixel<514) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=514 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=519 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=524 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=539 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=555 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=560 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=582 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=593 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=595 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=611 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=625 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=377 && xPixel<378 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=13 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=15 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=17 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=63 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=65 && yPixel<79) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=79 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=90 && yPixel<96) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=99 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=100 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=104 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=108 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=125 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=138 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=149 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=166 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=201 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=204 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=216 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=219 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=227 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=234 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=244 && yPixel<249) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=249 && yPixel<258) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=258 && yPixel<268) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=268 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=308 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=316 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=319 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=323 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=331 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=350 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=359 && yPixel<360) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=361 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=380 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=387 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=390 && yPixel<407) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=407 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=445 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=453 && yPixel<466) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=466 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=512 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=517 && yPixel<519) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=519 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=526 && yPixel<528) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=528 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=536 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=542 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=545 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=548 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=558 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=559 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=567 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=578 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=592 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=601 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=609 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=378 && xPixel<379 && yPixel>=617 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=13 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=36 && yPixel<45) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=47 && yPixel<51) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=51 && yPixel<54) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=55 && yPixel<59) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=59 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=64 && yPixel<76) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=76 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=86 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=89 && yPixel<98) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=98 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=106 && yPixel<111) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=111 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=123 && yPixel<125) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=125 && yPixel<127) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=127 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=134 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=136 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=141 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=146 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=150 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=163 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=187 && yPixel<190) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=190 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=195 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=203 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=211 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=225 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=231 && yPixel<235) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=237 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=240 && yPixel<244) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=244 && yPixel<247) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=247 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=250 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=253 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=257 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=266 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=268 && yPixel<278) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=278 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=321 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=327 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=332 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=338 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=341 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=349 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=366 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=369 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=385 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=400 && yPixel<405) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=405 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=416 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=437 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=445 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=483 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=501 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=516 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=522 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=527 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=534 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=536 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=557 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=571 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=587 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=603 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=608 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=612 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=379 && xPixel<380 && yPixel>=616 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=0 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=4 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=51 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=59 && yPixel<79) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=79 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=100 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=101 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=102 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=115 && yPixel<116) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=116 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=126 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=128 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=136 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=141 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=154 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=158 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=167 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=171 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=190 && yPixel<194) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=195 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=215 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=227 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=230 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=239 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=246 && yPixel<254) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=254 && yPixel<256) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=256 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=265 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=269 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=273 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=274 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=279 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=285 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=300 && yPixel<304) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=304 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=321 && yPixel<329) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=337 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=342 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=354 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=356 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=362 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=394 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=408 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=437 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=445 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=455 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=456 && yPixel<466) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=466 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=495 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=506 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=511 && yPixel<514) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=514 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=517 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=527 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=532 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=547 && yPixel<557) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=557 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=563 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=564 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=574 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=582 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=589 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=601 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=608 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=618 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=380 && xPixel<381 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=21 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=27 && yPixel<36) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=39 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=45 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=49 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=51 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=59 && yPixel<76) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=76 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=78 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=90 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=96 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=98 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=106 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=141 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=152 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=161 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=172 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=196 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=202 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=220 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=224 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=235 && yPixel<242) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=242 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=246 && yPixel<252) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=252 && yPixel<255) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=255 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=266 && yPixel<267) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=267 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=275 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=277 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=280 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=287 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=300 && yPixel<302) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=302 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=339 && yPixel<341) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=341 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=342 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=350 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=364 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=381 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=385 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=402 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=419 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=428 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=437 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=452 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=459 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=461 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=463 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=495 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=500 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=521 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=526 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=527 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=537 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=565 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=569 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=570 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=582 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=589 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=597 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=608 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=612 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=617 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=619 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=625 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=632 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=634 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=381 && xPixel<382 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=0 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=30 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=34 && yPixel<72) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=72 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=93 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=96 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=97 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=99 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=107 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=110 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=132 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=144 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=147 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=150 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=154 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=161 && yPixel<165) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=167 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=170 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=177 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=192 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=196 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=207 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=219 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=223 && yPixel<231) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=232 && yPixel<251) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=251 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=261 && yPixel<266) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=269 && yPixel<275) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=275 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=283 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=292 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=295 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=298 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=299 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=305 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=322 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=326 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=329 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=343 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=353 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=360 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=374 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=383 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=394 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=399 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=419 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=427 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=430 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=434 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=437 && yPixel<443) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=447 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=454 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=456 && yPixel<471) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=471 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=490 && yPixel<493) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=493 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=494 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=504 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=505 && yPixel<537) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=539 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=546 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=559 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=563 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=568 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=569 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=572 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=573 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=584 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=588 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=592 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=596 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=598 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=607 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=611 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=612 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=616 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=621 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=382 && xPixel<383 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=0 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=5 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=36 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=41 && yPixel<58) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=58 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=76 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=83 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=103 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=105 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=108 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=140 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=157 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=160 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=164 && yPixel<168) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=171 && yPixel<176) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=180 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=190 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=203 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=211 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=215 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=225 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=228 && yPixel<245) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=245 && yPixel<248) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=248 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=253 && yPixel<254) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=254 && yPixel<267) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=267 && yPixel<268) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=268 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=280 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=282 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=285 && yPixel<295) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=295 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=299 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=300 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=310 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=328 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=335 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=345 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=352 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=356 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=360 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=362 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=367 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=371 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=376 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=378 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=384 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=389 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=394 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=399 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=404 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=407 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=423 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=429 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=433 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=434 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=435 && yPixel<436) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=436 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=437 && yPixel<443) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=444 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=448 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=449 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=456 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=459 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=470 && yPixel<471) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=471 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=475 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=482 && yPixel<489) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=489 && yPixel<490) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=490 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=499 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=516 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=526 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=559 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=575 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=586 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=597 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=606 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=610 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=619 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=631 && yPixel<632) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=634 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=383 && xPixel<384 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=0 && yPixel<10) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=14 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=18 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=41 && yPixel<48) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=48 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=53 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=63 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=65 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=72 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=85 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=96 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=146 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=158 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=161 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=169 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=172 && yPixel<176) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=178 && yPixel<180) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=180 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=194 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=201 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=204 && yPixel<212) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=212 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=216 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=223 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=228 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=240 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=252 && yPixel<258) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=258 && yPixel<299) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=306 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=310 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=314 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=321 && yPixel<322) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=322 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=327 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=334 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=346 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=360 && yPixel<365) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=366 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=368 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=376 && yPixel<382) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=382 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=383 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=386 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=388 && yPixel<390) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=390 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=398 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=399 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=430 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=437 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=445 && yPixel<456) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=456 && yPixel<457) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=457 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=459 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=462 && yPixel<480) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=480 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=483 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=487 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=498 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=503 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=504 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=507 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=522 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=526 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=529 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=532 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=533 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=539 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=543 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=554 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=555 && yPixel<556) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=556 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=565 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=597 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=600 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=605 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=384 && xPixel<385 && yPixel>=606 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=20 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=38 && yPixel<47) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=50 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=52 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=55 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=56 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=79 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=83 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=99 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=107 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=114 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=144 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=158 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=168 && yPixel<180) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=182 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=185 && yPixel<186) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=186 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=194 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=208 && yPixel<214) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=217 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=233 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=263 && yPixel<277) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=277 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=279 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=297 && yPixel<301) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=301 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=303 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=308 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=323 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=327 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=335 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=344 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=355 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=361 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=365 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=367 && yPixel<379) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=383 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=384 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=391 && yPixel<401) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=401 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=404 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=405 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=409 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=411 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=446 && yPixel<449) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=449 && yPixel<454) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=454 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=475 && yPixel<482) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=482 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=483 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=490 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=494 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=498 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=505 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=509 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=528 && yPixel<529) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=529 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=536 && yPixel<543) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=546 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b11000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=562 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=565 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=566 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=577 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=581 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=585 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=596 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=385 && xPixel<386 && yPixel>=619 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=18 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=22 && yPixel<26) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=27 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=38 && yPixel<45) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=46 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=60 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=61 && yPixel<65) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=65 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=72 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=82 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=88 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=93 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=114 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=122 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=129 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=132 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b10000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=146 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=155 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=157 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=167 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=173 && yPixel<175) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=176 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=178 && yPixel<179) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=180 && yPixel<182) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=182 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=184 && yPixel<187) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=187 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=193 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=207 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=227 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=241 && yPixel<258) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=258 && yPixel<276) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=276 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=289 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=311 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=312 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=315 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=323 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=326 && yPixel<330) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=330 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=333 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=337 && yPixel<340) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=340 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=344 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=360 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=372 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=379 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=387 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=390 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=391 && yPixel<403) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=403 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=408 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=416 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=445 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=454 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=455 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=460 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=464 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=473 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=486 && yPixel<499) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=499 && yPixel<508) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=508 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=516 && yPixel<518) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=518 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=538 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=539 && yPixel<544) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=544 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=548 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=552 && yPixel<564) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=564 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=570 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=579 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=590 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=601 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=606 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=620 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=386 && xPixel<387 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=0 && yPixel<20) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=20 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=39 && yPixel<44) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=45 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=54 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=66 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=71 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=77 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=79 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=83 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=87 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=90 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=99 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=103 && yPixel<111) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=111 && yPixel<119) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=119 && yPixel<121) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=124 && yPixel<125) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=125 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=129 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=145 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=174 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=182 && yPixel<185) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=185 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=189 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=191 && yPixel<195) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=195 && yPixel<200) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=200 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=212 && yPixel<218) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=218 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=231 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=251 && yPixel<258) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=258 && yPixel<277) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=277 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=292 && yPixel<295) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=295 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=310 && yPixel<313) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=313 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=314 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=318 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=346 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=356 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=385 && yPixel<393) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=393 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=394 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=407 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=416 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=421 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=438 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=445 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=465 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=468 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=473 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=516 && yPixel<518) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=518 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=522 && yPixel<533) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=533 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=540 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=552 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=553 && yPixel<555) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=555 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=563 && yPixel<569) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=569 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=573 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=576 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=587 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=602 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=610 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=618 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=387 && xPixel<388 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=8 && yPixel<10) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=10 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=11 && yPixel<20) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=20 && yPixel<26) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=29 && yPixel<38) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=39 && yPixel<48) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=49 && yPixel<53) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=53 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=98 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=102 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=107 && yPixel<116) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=116 && yPixel<127) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=127 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=137 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=145 && yPixel<172) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=172 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=181 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=189 && yPixel<191) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=193 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=202 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=208 && yPixel<211) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=211 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=217 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=227 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=232 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=246 && yPixel<281) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=281 && yPixel<294) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=294 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=309 && yPixel<310) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=310 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=315 && yPixel<317) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=317 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=320 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=327 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=330 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=392 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=394 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=395 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=403 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=410 && yPixel<421) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=421 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=423 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=439 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=453 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=470 && yPixel<473) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=473 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=478 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=487 && yPixel<491) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=491 && yPixel<498) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=498 && yPixel<503) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=503 && yPixel<517) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=517 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=520 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=526 && yPixel<534) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=534 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=550 && yPixel<560) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=560 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=568 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=573 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=584 && yPixel<586) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=586 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=589 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=600 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=607 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=618 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=625 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=626 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=629 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=631 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=388 && xPixel<389 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=0 && yPixel<7) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=7 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=16 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=30 && yPixel<38) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=38 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=44 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=52 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=58 && yPixel<66) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=66 && yPixel<68) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=70 && yPixel<72) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=72 && yPixel<103) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=103 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=106 && yPixel<120) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=120 && yPixel<121) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=122 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=132 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=143 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=151 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=166 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=173 && yPixel<181) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=182 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=188 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=197 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=224 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=229 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=247 && yPixel<283) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=283 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=294 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=295 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=297 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=303 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=312 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=318 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=323 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=356 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=363 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=372 && yPixel<375) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=375 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=387 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=403 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=432 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=439 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=445 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=451 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=452 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=463 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=486 && yPixel<487) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=487 && yPixel<494) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=494 && yPixel<500) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=500 && yPixel<505) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=505 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=511 && yPixel<516) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=516 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=520 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=526 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=530 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=536 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=540 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=545 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=553 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=577 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=602 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=608 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=622 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=629 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=389 && xPixel<390 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=0 && yPixel<8) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=8 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=15 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=23 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=27 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=34 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=35 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=53 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=91 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=96 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=104 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=105 && yPixel<111) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=111 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=132 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=134 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=135 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=145 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=147 && yPixel<150) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=153 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=158 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=167 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=202 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=210 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=222 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=226 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=229 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=247 && yPixel<262) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=262 && yPixel<287) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=287 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=294 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=302 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=307 && yPixel<324) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=326 && yPixel<333) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=333 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=337 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=343 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=349 && yPixel<354) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=354 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=368 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=372 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=400 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=410 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=420 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=424 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=433 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=435 && yPixel<438) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=439 && yPixel<443) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=444 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=474 && yPixel<492) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=492 && yPixel<499) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=499 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=500 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=523 && yPixel<535) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=535 && yPixel<536) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=536 && yPixel<539) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=539 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=541 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=546 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=558 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=573 && yPixel<580) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=580 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=583 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=598 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=602 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=611 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=630 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=390 && xPixel<391 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=0 && yPixel<15) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=16 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=18 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=43 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=46 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=62 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=101 && yPixel<103) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=103 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=113 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=133 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=136 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=147 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=149 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=158 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=168 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=211 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=217 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=225 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=231 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=254 && yPixel<259) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=259 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=268 && yPixel<269) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=272 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=273 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=285 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=290 && yPixel<311) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=313 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=315 && yPixel<316) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=316 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=324 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=327 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=332 && yPixel<336) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=336 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=349 && yPixel<352) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=352 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=354 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=362 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=374 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=404 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=411 && yPixel<430) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=430 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=432 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=433 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=439 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=444 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=486 && yPixel<494) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=494 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=505 && yPixel<506) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=506 && yPixel<509) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=509 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=511 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=531 && yPixel<533) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=533 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=540 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=546 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=547 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=550 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=553 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=560 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=565 && yPixel<583) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=586 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=589 && yPixel<590) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=590 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=595 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=600 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=612 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=617 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=391 && xPixel<392 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=0 && yPixel<9) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=9 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=19 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=23 && yPixel<67) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=67 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=68 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=72 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=91 && yPixel<94) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=95 && yPixel<110) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=110 && yPixel<114) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=114 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=130 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=136 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=141 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=155 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=161 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=166 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=172 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=179 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=197 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=207 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=216 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=221 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=231 && yPixel<272) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=272 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=281 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=283 && yPixel<290) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=290 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=291 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=326 && yPixel<328) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=331 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=342 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=357 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=362 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=373 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=388 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=401 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=411 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=412 && yPixel<431) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=431 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=432 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=439 && yPixel<444) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=445 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=453 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=487 && yPixel<498) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=498 && yPixel<506) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=506 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=507 && yPixel<540) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=540 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=541 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=545 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=551 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=554 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=559 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=566 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=569 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=571 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=575 && yPixel<586) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=587 && yPixel<594) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=594 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=598 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=606 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=613 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=616 && yPixel<617) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=619 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=631 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=392 && xPixel<393 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=7 && yPixel<8) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=9 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=19 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=26 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=45 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=53 && yPixel<56) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=56 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=58 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=68 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=72 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=79 && yPixel<80) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=80 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=84 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=90 && yPixel<101) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=101 && yPixel<105) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=105 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=110 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=142 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=154 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=162 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=176 && yPixel<181) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=182 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=185 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=206 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=212 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=216 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=219 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=245 && yPixel<253) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=253 && yPixel<257) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=257 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=274 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=278 && yPixel<283) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=284 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=299 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=304 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=306 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=308 && yPixel<312) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=312 && yPixel<314) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=314 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=318 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=346 && yPixel<350) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=350 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=359 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=361 && yPixel<362) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=362 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=368 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=389 && yPixel<400) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=402 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=405 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=406 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=407 && yPixel<408) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=408 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=410 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=418 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=432 && yPixel<434) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=434 && yPixel<439) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=439 && yPixel<440) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=440 && yPixel<442) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=447 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=455 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=461 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=462 && yPixel<482) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=482 && yPixel<505) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=505 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=511 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=512 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=520 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=524 && yPixel<527) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=527 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=531 && yPixel<559) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=559 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=561 && yPixel<562) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=562 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=572 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=600 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=603 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=607 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=610 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=612 && yPixel<620) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=620 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=623 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=627 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=393 && xPixel<394 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=2 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=6 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=15 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=16 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=44 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=45 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=50 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=51 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=52 && yPixel<54) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=54 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=55 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=63 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=76 && yPixel<80) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=80 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=102 && yPixel<107) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=107 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=108 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=109 && yPixel<111) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=111 && yPixel<127) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=127 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=132 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=139 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=142 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=155 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=173 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=180 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=195 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=199 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=202 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=216 && yPixel<237) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=237 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=244 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=250 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=252 && yPixel<265) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=265 && yPixel<266) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=266 && yPixel<269) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=269 && yPixel<272) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=276 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=279 && yPixel<286) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=286 && yPixel<292) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=292 && yPixel<305) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=305 && yPixel<326) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=326 && yPixel<349) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=349 && yPixel<353) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=353 && yPixel<356) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=356 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=357 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=361 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=363 && yPixel<367) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=367 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=370 && yPixel<387) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=387 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=399 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=404 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=409 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=411 && yPixel<420) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=420 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=426 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=442 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=444 && yPixel<452) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=452 && yPixel<460) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=460 && yPixel<463) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=463 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=467 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=472 && yPixel<484) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=484 && yPixel<510) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=510 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=521 && yPixel<529) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=529 && yPixel<549) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=549 && yPixel<553) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=553 && yPixel<561) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=561 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=563 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=572 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=576 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=592 && yPixel<594) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=594 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=596 && yPixel<601) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=601 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=603 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=611 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=613 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=627 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=394 && xPixel<395 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=1 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=2 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=29 && yPixel<51) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=51 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=68 && yPixel<69) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=69 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=90 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=95 && yPixel<96) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=96 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=102 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=108 && yPixel<111) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=111 && yPixel<121) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=121 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=122 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=129 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b10000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=134 && yPixel<136) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b10000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b10000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=138 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=144 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=148 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=164 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=166 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=174 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=180 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=193 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=195 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=198 && yPixel<201) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=201 && yPixel<216) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=216 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=227 && yPixel<234) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=234 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=249 && yPixel<273) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=273 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=338 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=345 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=360 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=364 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=366 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=384 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=388 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=389 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=411 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=420 && yPixel<422) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=422 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=432 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=443 && yPixel<444) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=444 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=453 && yPixel<455) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=455 && yPixel<461) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=461 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=470 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=472 && yPixel<476) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=476 && yPixel<477) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=477 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=525 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=531 && yPixel<532) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=532 && yPixel<542) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=542 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=576 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=578 && yPixel<593) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=593 && yPixel<596) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=596 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b11000000,8'b10000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=600 && yPixel<606) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=606 && yPixel<608) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=614 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=619 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=630 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=395 && xPixel<396 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=6 && yPixel<7) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=7 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=11 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=13 && yPixel<14) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=14 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=41 && yPixel<46) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=48 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=50 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=57 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=61 && yPixel<67) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=67 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=74 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=75 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=76 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=89 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=109 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=123 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b10000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=132 && yPixel<135) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=136 && yPixel<142) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=142 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=165 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=174 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=181 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=197 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=200 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=213 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=215 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=223 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=230 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=237 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=239 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=243 && yPixel<254) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=254 && yPixel<284) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=284 && yPixel<308) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=308 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=319 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=327 && yPixel<337) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=337 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=338 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=353 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=357 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=367 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=368 && yPixel<392) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=392 && yPixel<397) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=397 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=411 && yPixel<422) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=422 && yPixel<428) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=428 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=433 && yPixel<435) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=435 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=437 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=445 && yPixel<466) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=466 && yPixel<467) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=467 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=470 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=478 && yPixel<481) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=481 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=498 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=504 && yPixel<523) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=523 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=524 && yPixel<526) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=526 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=535 && yPixel<539) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=539 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=551 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=558 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=572 && yPixel<575) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=578 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=581 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=582 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=592 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=597 && yPixel<605) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=616 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=621 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=623 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=630 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=396 && xPixel<397 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=0 && yPixel<2) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=2 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=4 && yPixel<13) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=13 && yPixel<17) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=18 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=23 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=29 && yPixel<35) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=36 && yPixel<40) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=40 && yPixel<46) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=46 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=52 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=53 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=62 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=71 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=74 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=77 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=85 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=94 && yPixel<97) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=97 && yPixel<98) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=98 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=101 && yPixel<112) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=112 && yPixel<113) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=113 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=114 && yPixel<121) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=121 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=130 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=133 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=138 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=163 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=164 && yPixel<168) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=168 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=177 && yPixel<188) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=188 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=190 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=194 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=199 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=217 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=225 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=229 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=239 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=244 && yPixel<245) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=245 && yPixel<246) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=246 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=258 && yPixel<282) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=284 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=306 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=319 && yPixel<326) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=326 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=331 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=338 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=342 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=343 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=349 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=374 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=383 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=394 && yPixel<395) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=395 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=404 && yPixel<429) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=429 && yPixel<430) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=430 && yPixel<432) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=432 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=446 && yPixel<473) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=473 && yPixel<474) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=474 && yPixel<485) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=485 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=487 && yPixel<495) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=495 && yPixel<497) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=497 && yPixel<498) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=498 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=503 && yPixel<511) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=511 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=521 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=531 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=536 && yPixel<553) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=553 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=560 && yPixel<562) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=562 && yPixel<571) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=571 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=576 && yPixel<581) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=581 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=583 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=590 && yPixel<593) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=593 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=603 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=616 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=630 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=636 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=397 && xPixel<398 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=0 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=6 && yPixel<8) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=8 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=9 && yPixel<13) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=13 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=20 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=34 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=53 && yPixel<80) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=80 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=87 && yPixel<121) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=121 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=123 && yPixel<124) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=124 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=138 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=141 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=163 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=167 && yPixel<173) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=173 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=195 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=200 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=219 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=227 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=241 && yPixel<244) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=244 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=249 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=259 && yPixel<261) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=261 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=306 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=316 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=318 && yPixel<326) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=326 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=332 && yPixel<342) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=342 && yPixel<346) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=346 && yPixel<349) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=350 && yPixel<361) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=361 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=373 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=379 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=384 && yPixel<399) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=399 && yPixel<428) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=428 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=446 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=456 && yPixel<476) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=476 && yPixel<519) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=519 && yPixel<520) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=522 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=525 && yPixel<529) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=529 && yPixel<530) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=530 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=531 && yPixel<536) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=536 && yPixel<557) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=557 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=564 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=565 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=571 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=577 && yPixel<579) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=579 && yPixel<582) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=582 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=587 && yPixel<595) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=602 && yPixel<604) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=604 && yPixel<609) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=610 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=616 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=398 && xPixel<399 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=11 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=16 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=25 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=52 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=60 && yPixel<71) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=74 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=83 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=89 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=130 && yPixel<131) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=131 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=136 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=140 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=142 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=145 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=163 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=167 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=174 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=179 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=190 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=204 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=205 && yPixel<208) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=210 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=217 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=229 && yPixel<239) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=239 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=241 && yPixel<247) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=247 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=274 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=284 && yPixel<307) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=307 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=314 && yPixel<315) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=315 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=322 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=327 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=331 && yPixel<347) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=347 && yPixel<349) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=349 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=351 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=353 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=373 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=376 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=394 && yPixel<527) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=527 && yPixel<535) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=535 && yPixel<564) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=564 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=571 && yPixel<584) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=584 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=587 && yPixel<597) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=597 && yPixel<606) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=606 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=607 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=614 && yPixel<616) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=619 && yPixel<620) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=620 && yPixel<622) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=624 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=399 && xPixel<400 && yPixel>=633 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=11 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=15 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=42 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=50 && yPixel<62) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=62 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=77 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=83 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=84 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=88 && yPixel<100) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=100 && yPixel<108) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=108 && yPixel<116) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=116 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=117 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=132 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b10000000,8'b10000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b10000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=140 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=147 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=156 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=158 && yPixel<161) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=161 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=166 && yPixel<173) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=173 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=190 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=198 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=203 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=207 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=210 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=228 && yPixel<245) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=245 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=270 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=274 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=276 && yPixel<278) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=278 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=280 && yPixel<281) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=282 && yPixel<283) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=283 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=284 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=285 && yPixel<318) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=318 && yPixel<321) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=321 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=323 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=331 && yPixel<340) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=340 && yPixel<348) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=348 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=355 && yPixel<357) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=357 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=360 && yPixel<363) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=363 && yPixel<364) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=364 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=365 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=371 && yPixel<402) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=402 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=413 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=442 && yPixel<471) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=471 && yPixel<472) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=472 && yPixel<524) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=524 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=534 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=537 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=543 && yPixel<572) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=577 && yPixel<578) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=578 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=583 && yPixel<599) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=599 && yPixel<608) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=608 && yPixel<619) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=619 && yPixel<627) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=627 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=628 && yPixel<635) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=400 && xPixel<401 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=11 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=28 && yPixel<40) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=42 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=46 && yPixel<47) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=47 && yPixel<48) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=48 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=49 && yPixel<51) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=51 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=61 && yPixel<72) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=73 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=82 && yPixel<87) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=87 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=90 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=94 && yPixel<95) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=95 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=114 && yPixel<117) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=117 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=132 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=145 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=153 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=156 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=161 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=171 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=172 && yPixel<175) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=175 && yPixel<178) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=178 && yPixel<187) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=187 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=198 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=201 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=209 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=211 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=215 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=220 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=227 && yPixel<230) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=231 && yPixel<252) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=252 && yPixel<253) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=253 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=261 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=263 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=269 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=271 && yPixel<272) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=272 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=284 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=293 && yPixel<304) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=304 && yPixel<315) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=315 && yPixel<318) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=318 && yPixel<319) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=319 && yPixel<320) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=320 && yPixel<323) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=323 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=329 && yPixel<331) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=332 && yPixel<334) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=334 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=339 && yPixel<342) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=342 && yPixel<373) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=373 && yPixel<388) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=388 && yPixel<391) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=391 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=403 && yPixel<410) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=410 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=425 && yPixel<437) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=438 && yPixel<440) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=440 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=444 && yPixel<452) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=452 && yPixel<458) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=458 && yPixel<525) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=525 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=534 && yPixel<538) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=538 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=540 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=548 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=554 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=564 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=568 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=610 && yPixel<618) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=618 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=624 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=628 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=631 && yPixel<638) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=401 && xPixel<402 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=0 && yPixel<32) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=34 && yPixel<35) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=40 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=43 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=44 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=49 && yPixel<52) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=52 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=61 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=74 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=78 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=84 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=85 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=89 && yPixel<90) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=90 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=92 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=141 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=154 && yPixel<156) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=156 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=161 && yPixel<163) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=166 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=171 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=174 && yPixel<177) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=179 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=199 && yPixel<205) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=205 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=219 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=224 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=234 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=238 && yPixel<251) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=251 && yPixel<252) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=252 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=256 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=260 && yPixel<279) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=279 && yPixel<290) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=290 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=298 && yPixel<319) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=319 && yPixel<321) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=321 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=334 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=339 && yPixel<364) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=364 && yPixel<368) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=368 && yPixel<384) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=384 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=386 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=402 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=411 && yPixel<414) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=414 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=419 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=425 && yPixel<426) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=426 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=429 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=441 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=446 && yPixel<453) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=453 && yPixel<456) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=456 && yPixel<537) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=537 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=544 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=551 && yPixel<552) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=552 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=561 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=567 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=572 && yPixel<590) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=590 && yPixel<607) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=607 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=625 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=402 && xPixel<403 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=28 && yPixel<33) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=34 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=36 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=45 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=62 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=71 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=130 && yPixel<137) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=137 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=139 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=153 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=158 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=161 && yPixel<164) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=164 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=181 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=190 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=211 && yPixel<216) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=218 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=222 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=225 && yPixel<228) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=238 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=241 && yPixel<244) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=246 && yPixel<253) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=253 && yPixel<255) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=255 && yPixel<259) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=261 && yPixel<283) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=283 && yPixel<285) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=285 && yPixel<287) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=287 && yPixel<288) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=291 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=299 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=304 && yPixel<310) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=310 && yPixel<320) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=320 && yPixel<330) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=335 && yPixel<347) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=347 && yPixel<356) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=356 && yPixel<363) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=363 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=366 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=375 && yPixel<393) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=393 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=400 && yPixel<413) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=413 && yPixel<421) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=421 && yPixel<427) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=427 && yPixel<429) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=431 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=445 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=453 && yPixel<538) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=538 && yPixel<573) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=573 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=574 && yPixel<576) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=577 && yPixel<581) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=581 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=587 && yPixel<600) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=600 && yPixel<612) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=612 && yPixel<616) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=616 && yPixel<628) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=628 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=629 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=630 && yPixel<632) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=632 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=633 && yPixel<636) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=403 && xPixel<404 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=21 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=28 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=40 && yPixel<59) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=59 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=61 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=64 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=65 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=114 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=115 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=139 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=146 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=151 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=157 && yPixel<158) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=158 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=162 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=166 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=177 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=180 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=191 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=206 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=221 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=235 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=242 && yPixel<245) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=245 && yPixel<247) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=248 && yPixel<257) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=259 && yPixel<262) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=262 && yPixel<263) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=263 && yPixel<264) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=264 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=265 && yPixel<288) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=288 && yPixel<293) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=293 && yPixel<300) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=300 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=311 && yPixel<321) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=321 && yPixel<328) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=328 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=336 && yPixel<338) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=338 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=351 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=354 && yPixel<390) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=390 && yPixel<394) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=394 && yPixel<399) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=399 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=400 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=407 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=412 && yPixel<425) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=425 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=432 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=437 && yPixel<438) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=438 && yPixel<439) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=439 && yPixel<441) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=441 && yPixel<442) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=442 && yPixel<443) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=443 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=445 && yPixel<447) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=447 && yPixel<449) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=449 && yPixel<450) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=450 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=451 && yPixel<469) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=469 && yPixel<479) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=479 && yPixel<494) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=494 && yPixel<531) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=531 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=554 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=560 && yPixel<568) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=568 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=592 && yPixel<595) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=595 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=597 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=598 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=607 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=609 && yPixel<615) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=615 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=633 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=404 && xPixel<405 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=14 && yPixel<16) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=16 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=18 && yPixel<21) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=23 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=25 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=33 && yPixel<44) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=44 && yPixel<47) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=47 && yPixel<53) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=53 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=71 && yPixel<72) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=72 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=74 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=94 && yPixel<104) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=104 && yPixel<112) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=112 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=115 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=135 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=143 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=153 && yPixel<155) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=155 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=160 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=169 && yPixel<171) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=171 && yPixel<175) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=175 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=199 && yPixel<206) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=208 && yPixel<209) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=210 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=220 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=226 && yPixel<244) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=244 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=266 && yPixel<284) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=284 && yPixel<290) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=290 && yPixel<292) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=292 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=293 && yPixel<294) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=294 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=298 && yPixel<306) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=306 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=309 && yPixel<311) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=311 && yPixel<314) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=314 && yPixel<319) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=319 && yPixel<326) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=326 && yPixel<327) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=327 && yPixel<332) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=332 && yPixel<333) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=333 && yPixel<355) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=355 && yPixel<365) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=365 && yPixel<370) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=370 && yPixel<381) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=381 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=385 && yPixel<389) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=389 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=392 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=445 && yPixel<454) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=454 && yPixel<459) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=459 && yPixel<460) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=460 && yPixel<501) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=501 && yPixel<545) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=545 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=561 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=567 && yPixel<577) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=577 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=607 && yPixel<615) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=615 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=621 && yPixel<626) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=626 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=405 && xPixel<406 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=18 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=20 && yPixel<25) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=26 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=45 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=110 && yPixel<113) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=113 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=135 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=154 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=160 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=163 && yPixel<174) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=174 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=200 && yPixel<228) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=228 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=231 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=238 && yPixel<239) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=239 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=244 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=255 && yPixel<284) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=284 && yPixel<292) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=292 && yPixel<294) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=294 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=297 && yPixel<303) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=303 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=304 && yPixel<307) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=307 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=311 && yPixel<316) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=316 && yPixel<323) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=323 && yPixel<330) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=330 && yPixel<334) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=334 && yPixel<338) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=338 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=339 && yPixel<352) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=352 && yPixel<362) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=362 && yPixel<370) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=370 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=374 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=375 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=378 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=385 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=387 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=388 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=402 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=411 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=415 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=423 && yPixel<428) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=428 && yPixel<503) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=503 && yPixel<573) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=573 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=577 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=582 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=624 && yPixel<637) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=406 && xPixel<407 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=0 && yPixel<14) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=14 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=18 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=24 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=43 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=102 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=106 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=136 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=152 && yPixel<175) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=175 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=181 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=192 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=200 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=202 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=206 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=215 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=223 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=231 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=234 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=247 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=266 && yPixel<288) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=288 && yPixel<291) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=291 && yPixel<294) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=294 && yPixel<314) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=314 && yPixel<340) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=340 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=345 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=352 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=369 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=376 && yPixel<394) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=394 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=396 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=414 && yPixel<420) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=420 && yPixel<441) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=441 && yPixel<444) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=446 && yPixel<468) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=468 && yPixel<470) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=470 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=511 && yPixel<590) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=590 && yPixel<609) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=610 && yPixel<618) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=618 && yPixel<635) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=407 && xPixel<408 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=0 && yPixel<21) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=22 && yPixel<33) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=35 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=43 && yPixel<99) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=99 && yPixel<101) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=101 && yPixel<119) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=119 && yPixel<120) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=120 && yPixel<133) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=133 && yPixel<134) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=134 && yPixel<139) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=139 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=145 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=154 && yPixel<161) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=161 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=169 && yPixel<173) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=174 && yPixel<176) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=176 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=180 && yPixel<194) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=194 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=207 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=218 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=221 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=226 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=237 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=238 && yPixel<243) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=243 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=244 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=246 && yPixel<255) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=255 && yPixel<284) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=284 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=286 && yPixel<297) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=297 && yPixel<340) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=340 && yPixel<343) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=343 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=344 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=351 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=356 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=371 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=376 && yPixel<398) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=398 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=400 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=417 && yPixel<419) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=419 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=445 && yPixel<446) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=446 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=447 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=448 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=472 && yPixel<490) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=490 && yPixel<491) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=491 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=521 && yPixel<582) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=582 && yPixel<585) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=585 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=586 && yPixel<598) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=598 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=600 && yPixel<603) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=604 && yPixel<605) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=605 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=610 && yPixel<617) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=617 && yPixel<621) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=621 && yPixel<625) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=625 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=408 && xPixel<409 && yPixel>=631 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=18 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=19 && yPixel<30) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=33 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=39 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=69 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=78 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=79 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=82 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=83 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=132 && yPixel<133) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=133 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=136 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=141 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=143 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=150 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=151 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=154 && yPixel<155) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=155 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=159 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=163 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=167 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=171 && yPixel<190) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=190 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=193 && yPixel<195) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=195 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=198 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=207 && yPixel<211) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=211 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=214 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=220 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=227 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=230 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=236 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=241 && yPixel<245) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=245 && yPixel<272) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=272 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=345 && yPixel<348) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=348 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=350 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=353 && yPixel<354) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=354 && yPixel<362) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=362 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=374 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=383 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=387 && yPixel<392) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=392 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=401 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=415 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=418 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=452 && yPixel<453) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=453 && yPixel<462) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=462 && yPixel<472) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=472 && yPixel<480) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=480 && yPixel<523) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=523 && yPixel<582) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=582 && yPixel<584) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=584 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=585 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=597 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=603 && yPixel<634) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=634 && yPixel<635) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=635 && yPixel<637) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=409 && xPixel<410 && yPixel>=637 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=3 && yPixel<4) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=4 && yPixel<5) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=5 && yPixel<6) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=6 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=19 && yPixel<20) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=20 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=21 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=22 && yPixel<23) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=23 && yPixel<24) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=24 && yPixel<30) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=30 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=33 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=38 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=65 && yPixel<75) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=75 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=77 && yPixel<84) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=84 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=92 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=94 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=108 && yPixel<113) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=113 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=115 && yPixel<120) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=120 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=122 && yPixel<125) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=125 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=131 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=136 && yPixel<137) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=137 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=147 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=148 && yPixel<149) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=149 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=156 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=164 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=166 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=170 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=176 && yPixel<192) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=192 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=210 && yPixel<211) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=214 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=218 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=221 && yPixel<225) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=226 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=233 && yPixel<234) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=234 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=241 && yPixel<256) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=256 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=259 && yPixel<281) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=281 && yPixel<282) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=282 && yPixel<298) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=298 && yPixel<308) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=308 && yPixel<311) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=311 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=313 && yPixel<332) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=332 && yPixel<342) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=342 && yPixel<345) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=345 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=346 && yPixel<351) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=351 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=359 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=375 && yPixel<376) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=376 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=377 && yPixel<385) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=385 && yPixel<409) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=409 && yPixel<457) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=457 && yPixel<464) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=464 && yPixel<470) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=470 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=477 && yPixel<481) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=481 && yPixel<486) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=486 && yPixel<491) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=491 && yPixel<525) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=525 && yPixel<589) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=589 && yPixel<594) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=595 && yPixel<598) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=598 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=599 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=600 && yPixel<601) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=601 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=602 && yPixel<603) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=603 && yPixel<610) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=610 && yPixel<611) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=611 && yPixel<616) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=616 && yPixel<624) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=624 && yPixel<636) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=410 && xPixel<411 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=0 && yPixel<1) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=1 && yPixel<3) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=3 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=18 && yPixel<21) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=21 && yPixel<28) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=33 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=39 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=41 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=46 && yPixel<57) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=57 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=58 && yPixel<62) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=62 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=64 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=71 && yPixel<77) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=77 && yPixel<78) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=78 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=81 && yPixel<83) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=83 && yPixel<85) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=85 && yPixel<86) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=86 && yPixel<92) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=92 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=94 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=108 && yPixel<112) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=112 && yPixel<115) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=115 && yPixel<117) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=117 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=141 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=151 && yPixel<152) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=153 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=160 && yPixel<170) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=170 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=173 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=177 && yPixel<181) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=181 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=194 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=198 && yPixel<201) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=201 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=207 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=210 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=213 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=221 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=223 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=230 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=232 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=233 && yPixel<265) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=265 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=270 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=274 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=297 && yPixel<312) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=312 && yPixel<313) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=313 && yPixel<325) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=325 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=329 && yPixel<334) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=334 && yPixel<358) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=358 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=359 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=369 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=370 && yPixel<372) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=372 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=377 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=401 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=403 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=413 && yPixel<416) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=416 && yPixel<472) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=472 && yPixel<475) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=475 && yPixel<477) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=477 && yPixel<478) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=478 && yPixel<483) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=483 && yPixel<489) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=489 && yPixel<528) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=528 && yPixel<590) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=590 && yPixel<596) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=596 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=599 && yPixel<627) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=627 && yPixel<636) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=411 && xPixel<412 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=3 && yPixel<5) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=5 && yPixel<9) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=9 && yPixel<15) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=15 && yPixel<25) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=25 && yPixel<28) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=29 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=33 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=43 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=46 && yPixel<55) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=55 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=58 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=65 && yPixel<83) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=83 && yPixel<88) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=88 && yPixel<89) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=89 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=92 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=140 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=143 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=154 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=160 && yPixel<165) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=168 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=175 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=177 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=178 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=199 && yPixel<208) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=208 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=210 && yPixel<212) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=212 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=217 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=220 && yPixel<222) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=222 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=223 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=225 && yPixel<229) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=231 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=243 && yPixel<246) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=246 && yPixel<247) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=247 && yPixel<248) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=248 && yPixel<306) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=306 && yPixel<324) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=324 && yPixel<328) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=328 && yPixel<331) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=332 && yPixel<342) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=342 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=347 && yPixel<358) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=358 && yPixel<360) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=360 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=369 && yPixel<371) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=371 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=376 && yPixel<403) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=403 && yPixel<404) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=404 && yPixel<413) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=413 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=415 && yPixel<445) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=445 && yPixel<448) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=448 && yPixel<450) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=450 && yPixel<462) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=462 && yPixel<477) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=477 && yPixel<500) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=500 && yPixel<517) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=517 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=526 && yPixel<573) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=573 && yPixel<575) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=575 && yPixel<576) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=577 && yPixel<610) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=610 && yPixel<615) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=615 && yPixel<616) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=616 && yPixel<619) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=621 && yPixel<632) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=412 && xPixel<413 && yPixel>=632 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=0 && yPixel<25) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=25 && yPixel<27) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=27 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=31 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=33 && yPixel<35) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=35 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=36 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=41 && yPixel<58) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=58 && yPixel<61) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=61 && yPixel<68) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=68 && yPixel<70) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=70 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=71 && yPixel<73) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=73 && yPixel<74) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=74 && yPixel<76) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=76 && yPixel<93) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=93 && yPixel<94) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=94 && yPixel<140) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=140 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=144 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=153 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=169 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=173 && yPixel<174) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=174 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=175 && yPixel<186) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=186 && yPixel<187) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=192 && yPixel<193) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=193 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=195 && yPixel<203) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=203 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=209 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=212 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=218 && yPixel<224) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=224 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=226 && yPixel<238) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=238 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=241 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=242 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=261 && yPixel<262) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=262 && yPixel<269) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=269 && yPixel<270) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=270 && yPixel<271) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=271 && yPixel<274) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=274 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=275 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=280 && yPixel<285) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=285 && yPixel<286) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=286 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=289 && yPixel<310) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=310 && yPixel<328) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=328 && yPixel<333) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=333 && yPixel<336) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=336 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=337 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=365 && yPixel<366) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=366 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=367 && yPixel<372) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=372 && yPixel<373) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=373 && yPixel<378) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=380 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=400 && yPixel<401) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=407 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=444 && yPixel<446) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=446 && yPixel<452) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=452 && yPixel<576) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=576 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=577 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=585 && yPixel<598) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=598 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=607 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=614 && yPixel<621) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=621 && yPixel<624) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=413 && xPixel<414 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=0 && yPixel<27) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=27 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=32 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=34 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=38 && yPixel<39) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=39 && yPixel<91) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=91 && yPixel<92) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=92 && yPixel<116) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=116 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=130 && yPixel<142) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=143 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=145 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=146 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=149 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=151 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=154 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=165 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=170 && yPixel<187) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=187 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=192 && yPixel<199) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=199 && yPixel<202) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=206 && yPixel<207) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=207 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=215 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=217 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=221 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=224 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=227 && yPixel<259) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=259 && yPixel<264) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=264 && yPixel<273) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=273 && yPixel<275) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=275 && yPixel<276) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=276 && yPixel<277) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=277 && yPixel<279) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=279 && yPixel<280) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=280 && yPixel<284) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=288 && yPixel<297) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=297 && yPixel<309) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=309 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=324 && yPixel<329) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=329 && yPixel<352) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=352 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=359 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=371 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=384 && yPixel<388) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=388 && yPixel<405) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=405 && yPixel<444) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=444 && yPixel<445) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=445 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=451 && yPixel<532) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=532 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=551 && yPixel<578) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=578 && yPixel<579) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=579 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=580 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=585 && yPixel<589) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=589 && yPixel<613) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=613 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=626 && yPixel<630) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=631 && yPixel<633) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=633 && yPixel<635) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=414 && xPixel<415 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=0 && yPixel<24) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=24 && yPixel<25) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=25 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=27 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=31 && yPixel<36) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=36 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=37 && yPixel<38) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=38 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=41 && yPixel<65) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=65 && yPixel<69) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=69 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=71 && yPixel<76) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=76 && yPixel<79) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=79 && yPixel<82) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=82 && yPixel<105) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=105 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=128 && yPixel<129) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=129 && yPixel<130) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=130 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=141 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=144 && yPixel<149) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=149 && yPixel<152) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=152 && yPixel<153) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=153 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=170 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=177 && yPixel<179) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=179 && yPixel<180) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=180 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=185 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=219 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=226 && yPixel<227) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=227 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=234 && yPixel<235) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=235 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=249 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=251 && yPixel<257) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=257 && yPixel<259) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=259 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=260 && yPixel<272) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=272 && yPixel<284) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=284 && yPixel<288) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=288 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=289 && yPixel<295) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=295 && yPixel<296) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=296 && yPixel<302) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=302 && yPixel<308) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=308 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=349 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=350 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=368 && yPixel<386) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=386 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=387 && yPixel<414) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=414 && yPixel<417) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=417 && yPixel<456) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=456 && yPixel<493) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=493 && yPixel<504) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=504 && yPixel<507) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=507 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=512 && yPixel<531) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=531 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=537 && yPixel<538) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=541 && yPixel<544) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=544 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=546 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=556 && yPixel<561) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=561 && yPixel<583) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=583 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=586 && yPixel<597) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=597 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=610 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=619 && yPixel<634) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=415 && xPixel<416 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=26 && yPixel<27) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=27 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=28 && yPixel<39) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=41 && yPixel<45) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=45 && yPixel<46) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=46 && yPixel<49) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=49 && yPixel<50) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=50 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=60 && yPixel<80) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=80 && yPixel<81) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=81 && yPixel<82) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=82 && yPixel<102) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=102 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=135 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=138 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=143 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=146 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=147 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=157 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=160 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=164 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=172 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=173 && yPixel<175) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=175 && yPixel<181) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=181 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=183 && yPixel<193) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=193 && yPixel<196) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=196 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=198 && yPixel<210) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=210 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=214 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=216 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=221 && yPixel<226) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=226 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=239 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=248 && yPixel<249) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=249 && yPixel<256) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=256 && yPixel<279) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=279 && yPixel<286) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=286 && yPixel<289) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=289 && yPixel<293) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=293 && yPixel<299) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=299 && yPixel<322) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=322 && yPixel<330) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=330 && yPixel<343) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=343 && yPixel<350) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=350 && yPixel<367) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=367 && yPixel<370) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=370 && yPixel<377) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=377 && yPixel<381) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=381 && yPixel<383) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=383 && yPixel<387) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=387 && yPixel<410) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=411 && yPixel<415) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=415 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=432 && yPixel<465) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=465 && yPixel<500) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=500 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=548 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=551 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=553 && yPixel<558) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=558 && yPixel<560) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=560 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=565 && yPixel<590) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=590 && yPixel<592) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=592 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=599 && yPixel<603) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=603 && yPixel<604) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=604 && yPixel<613) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=613 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=622 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=416 && xPixel<417 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=17 && yPixel<19) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=19 && yPixel<34) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=34 && yPixel<37) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=37 && yPixel<79) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=79 && yPixel<112) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=112 && yPixel<124) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=124 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=132 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=135 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=139 && yPixel<142) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=144 && yPixel<145) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=145 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=163 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=165 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=166 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=169 && yPixel<175) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=175 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=178 && yPixel<183) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=183 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=184 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=191 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=194 && yPixel<195) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=195 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=197 && yPixel<202) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=202 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=206 && yPixel<208) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=208 && yPixel<211) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=211 && yPixel<212) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=212 && yPixel<214) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=220 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=229 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=231 && yPixel<232) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=232 && yPixel<234) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=234 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=236 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=240 && yPixel<241) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=241 && yPixel<248) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=248 && yPixel<253) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=253 && yPixel<262) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=262 && yPixel<284) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=284 && yPixel<293) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=293 && yPixel<296) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=296 && yPixel<297) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=297 && yPixel<298) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=298 && yPixel<304) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=304 && yPixel<344) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=344 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=347 && yPixel<351) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=351 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=356 && yPixel<375) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=375 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=384 && yPixel<406) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=406 && yPixel<432) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=432 && yPixel<473) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=473 && yPixel<498) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=498 && yPixel<512) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=512 && yPixel<525) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=525 && yPixel<541) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=541 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=546 && yPixel<550) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=551 && yPixel<565) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=565 && yPixel<569) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=569 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=574 && yPixel<594) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=599 && yPixel<602) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=602 && yPixel<607) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=607 && yPixel<610) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=610 && yPixel<614) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=615 && yPixel<619) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=619 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=621 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=627 && yPixel<629) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=417 && xPixel<418 && yPixel>=629 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=0 && yPixel<17) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=17 && yPixel<18) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=18 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=39 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=40 && yPixel<73) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=73 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=106 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=110 && yPixel<114) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=114 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=132 && yPixel<136) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=138 && yPixel<147) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=147 && yPixel<151) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=151 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=154 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=163 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=166 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=168 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=170 && yPixel<184) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=184 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=191 && yPixel<200) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=200 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=216 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=217 && yPixel<219) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=220 && yPixel<223) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=223 && yPixel<224) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=227 && yPixel<228) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=228 && yPixel<229) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=229 && yPixel<230) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=230 && yPixel<231) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=231 && yPixel<235) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=235 && yPixel<236) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=236 && yPixel<237) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=237 && yPixel<247) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=247 && yPixel<256) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=256 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=260 && yPixel<266) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=266 && yPixel<290) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=290 && yPixel<296) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=296 && yPixel<299) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=299 && yPixel<301) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=301 && yPixel<305) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=305 && yPixel<318) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=318 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=327 && yPixel<346) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=346 && yPixel<353) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=353 && yPixel<355) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=355 && yPixel<356) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=356 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=368 && yPixel<369) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=369 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=371 && yPixel<376) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=376 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=382 && yPixel<384) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=384 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=423 && yPixel<424) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=424 && yPixel<447) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=447 && yPixel<451) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=451 && yPixel<465) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=465 && yPixel<468) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=468 && yPixel<480) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=480 && yPixel<495) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=495 && yPixel<537) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=537 && yPixel<543) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=543 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=546 && yPixel<563) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=563 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=577 && yPixel<598) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=598 && yPixel<608) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=608 && yPixel<609) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=609 && yPixel<612) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=612 && yPixel<621) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=621 && yPixel<622) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=622 && yPixel<623) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=623 && yPixel<626) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=626 && yPixel<627) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=627 && yPixel<630) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=630 && yPixel<631) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=631 && yPixel<636) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=418 && xPixel<419 && yPixel>=636 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=0 && yPixel<18) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=18 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=22 && yPixel<40) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=40 && yPixel<41) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=41 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=42 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=43 && yPixel<59) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=59 && yPixel<60) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=60 && yPixel<62) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=62 && yPixel<106) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=106 && yPixel<108) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=108 && yPixel<122) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=122 && yPixel<123) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=123 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=126 && yPixel<129) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=129 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=131 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=139 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=143 && yPixel<150) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=150 && yPixel<156) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=156 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=159 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=160 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=162 && yPixel<166) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=166 && yPixel<178) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=178 && yPixel<181) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=181 && yPixel<182) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=182 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=188 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=197 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=203 && yPixel<213) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=213 && yPixel<216) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=216 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=221 && yPixel<225) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=225 && yPixel<227) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=227 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=233 && yPixel<242) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=242 && yPixel<243) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=243 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=260 && yPixel<274) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=274 && yPixel<294) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=294 && yPixel<303) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=303 && yPixel<308) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=308 && yPixel<309) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=309 && yPixel<324) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=324 && yPixel<327) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=327 && yPixel<365) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=365 && yPixel<368) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=368 && yPixel<371) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=371 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=377 && yPixel<385) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=385 && yPixel<396) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=396 && yPixel<400) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=400 && yPixel<402) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=402 && yPixel<423) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=423 && yPixel<425) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=425 && yPixel<481) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=481 && yPixel<498) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=498 && yPixel<508) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=508 && yPixel<511) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=511 && yPixel<529) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=529 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=531 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=567 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=574 && yPixel<575) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=575 && yPixel<577) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=577 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=607 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=614 && yPixel<617) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=617 && yPixel<624) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=624 && yPixel<625) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=419 && xPixel<420 && yPixel>=625 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=0 && yPixel<29) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=29 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=33 && yPixel<39) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=39 && yPixel<43) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=43 && yPixel<55) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=55 && yPixel<69) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=69 && yPixel<71) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=71 && yPixel<126) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=126 && yPixel<128) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=128 && yPixel<132) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=132 && yPixel<137) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=137 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=142 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=144 && yPixel<146) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=146 && yPixel<148) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=148 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=151 && yPixel<157) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=157 && yPixel<159) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=159 && yPixel<161) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=162 && yPixel<163) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=163 && yPixel<170) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=170 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=171 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=176 && yPixel<182) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=182 && yPixel<185) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=185 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=188 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=200 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=203 && yPixel<204) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=204 && yPixel<212) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=212 && yPixel<213) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=213 && yPixel<214) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=214 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=220 && yPixel<221) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=221 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=239 && yPixel<240) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=240 && yPixel<242) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=242 && yPixel<258) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=258 && yPixel<260) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=260 && yPixel<261) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=261 && yPixel<268) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=268 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=280 && yPixel<304) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=304 && yPixel<313) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=313 && yPixel<316) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=316 && yPixel<348) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=348 && yPixel<359) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=359 && yPixel<374) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=374 && yPixel<377) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=377 && yPixel<382) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=382 && yPixel<386) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=386 && yPixel<412) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=412 && yPixel<418) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=418 && yPixel<427) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=427 && yPixel<433) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=433 && yPixel<486) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=486 && yPixel<498) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=498 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=507 && yPixel<509) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=509 && yPixel<513) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=513 && yPixel<517) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=517 && yPixel<527) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=527 && yPixel<531) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=531 && yPixel<545) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=545 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=546 && yPixel<548) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=548 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=550 && yPixel<554) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=554 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=567 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=570 && yPixel<573) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=573 && yPixel<580) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=580 && yPixel<582) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=582 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=583 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=614 && yPixel<618) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=619 && yPixel<624) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=420 && xPixel<421 && yPixel>=624 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=0 && yPixel<19) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=19 && yPixel<22) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=22 && yPixel<53) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=53 && yPixel<135) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=135 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=139 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=141 && yPixel<147) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=147 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=151 && yPixel<153) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=153 && yPixel<154) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=154 && yPixel<164) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=164 && yPixel<168) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=168 && yPixel<171) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=171 && yPixel<173) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=173 && yPixel<175) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=175 && yPixel<176) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=176 && yPixel<177) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=177 && yPixel<188) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=188 && yPixel<191) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=191 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=198 && yPixel<202) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=202 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=203 && yPixel<214) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=214 && yPixel<217) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=217 && yPixel<218) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=218 && yPixel<219) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=219 && yPixel<220) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=220 && yPixel<239) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=239 && yPixel<244) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=244 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=280 && yPixel<316) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=316 && yPixel<324) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=324 && yPixel<328) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=328 && yPixel<329) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=329 && yPixel<345) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=345 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=347 && yPixel<357) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=357 && yPixel<368) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=368 && yPixel<411) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=411 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=429 && yPixel<434) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=434 && yPixel<437) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=437 && yPixel<505) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=505 && yPixel<507) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=507 && yPixel<520) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=520 && yPixel<521) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=521 && yPixel<522) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=522 && yPixel<524) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=524 && yPixel<525) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=525 && yPixel<526) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=526 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=547 && yPixel<552) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=552 && yPixel<566) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=566 && yPixel<567) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=567 && yPixel<568) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=568 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=574 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=583 && yPixel<585) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=585 && yPixel<587) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=587 && yPixel<589) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=589 && yPixel<594) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=594 && yPixel<599) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=599 && yPixel<609) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=609 && yPixel<610) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=610 && yPixel<626) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=626 && yPixel<628) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=628 && yPixel<634) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=421 && xPixel<422 && yPixel>=634 && yPixel<639) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=0 && yPixel<3) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=3 && yPixel<12) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=12 && yPixel<13) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=13 && yPixel<23) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=23 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=28 && yPixel<30) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=30 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=33 && yPixel<34) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=34 && yPixel<42) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=42 && yPixel<51) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=51 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=136 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=146 && yPixel<161) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=161 && yPixel<162) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=162 && yPixel<167) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=167 && yPixel<168) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=168 && yPixel<169) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=169 && yPixel<170) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=170 && yPixel<172) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=172 && yPixel<186) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=186 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=191 && yPixel<193) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=193 && yPixel<198) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=199 && yPixel<200) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=200 && yPixel<201) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=201 && yPixel<204) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=204 && yPixel<207) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=207 && yPixel<209) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=209 && yPixel<210) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=210 && yPixel<215) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=215 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=217 && yPixel<233) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=233 && yPixel<241) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=241 && yPixel<251) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=251 && yPixel<256) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=256 && yPixel<280) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=280 && yPixel<300) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=300 && yPixel<307) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=307 && yPixel<312) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=312 && yPixel<327) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=327 && yPixel<331) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=331 && yPixel<335) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=335 && yPixel<337) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=337 && yPixel<347) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=347 && yPixel<349) {VGAr,VGAg,VRAb}={8'b11000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=349 && yPixel<353) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=353 && yPixel<360) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=360 && yPixel<379) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=379 && yPixel<406) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=406 && yPixel<410) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=410 && yPixel<411) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=411 && yPixel<416) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=418 && yPixel<420) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=420 && yPixel<436) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=436 && yPixel<487) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=487 && yPixel<503) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=503 && yPixel<513) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=513 && yPixel<534) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=534 && yPixel<538) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=538 && yPixel<541) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=541 && yPixel<546) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=546 && yPixel<563) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=563 && yPixel<565) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=565 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=574 && yPixel<583) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=583 && yPixel<584) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=584 && yPixel<588) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=588 && yPixel<607) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=607 && yPixel<612) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=612 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=614 && yPixel<615) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=615 && yPixel<618) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=618 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=623 && yPixel<635) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=422 && xPixel<423 && yPixel>=635 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=0 && yPixel<26) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=26 && yPixel<28) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=28 && yPixel<29) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=29 && yPixel<31) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=31 && yPixel<32) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=32 && yPixel<33) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=33 && yPixel<109) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=109 && yPixel<110) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=110 && yPixel<116) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=116 && yPixel<117) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=117 && yPixel<136) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=136 && yPixel<138) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=138 && yPixel<139) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=139 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=144 && yPixel<157) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=157 && yPixel<160) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=160 && yPixel<165) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=165 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=167 && yPixel<180) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=180 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=184 && yPixel<187) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=187 && yPixel<188) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=188 && yPixel<189) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=189 && yPixel<190) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=190 && yPixel<191) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=191 && yPixel<192) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=192 && yPixel<194) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=194 && yPixel<196) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=196 && yPixel<197) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=198 && yPixel<208) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=208 && yPixel<212) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=212 && yPixel<215) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=215 && yPixel<224) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=224 && yPixel<225) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=225 && yPixel<226) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=226 && yPixel<233) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=233 && yPixel<249) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=249 && yPixel<250) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=250 && yPixel<261) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=261 && yPixel<278) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=278 && yPixel<316) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=316 && yPixel<320) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=320 && yPixel<329) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=329 && yPixel<330) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=330 && yPixel<335) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=335 && yPixel<354) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=354 && yPixel<379) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=381 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=393 && yPixel<396) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=396 && yPixel<399) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=399 && yPixel<402) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=402 && yPixel<404) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=404 && yPixel<414) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=414 && yPixel<416) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=418 && yPixel<419) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=419 && yPixel<422) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=422 && yPixel<423) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=423 && yPixel<426) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=426 && yPixel<443) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=443 && yPixel<463) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=463 && yPixel<516) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=516 && yPixel<540) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=540 && yPixel<547) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=547 && yPixel<570) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=570 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11111111,8'b10000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=572 && yPixel<574) {VGAr,VGAg,VRAb}={8'b11111111,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=574 && yPixel<583) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=583 && yPixel<588) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=588 && yPixel<589) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=589 && yPixel<594) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=594 && yPixel<614) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=614 && yPixel<619) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=619 && yPixel<623) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=623 && yPixel<625) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=625 && yPixel<629) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=629 && yPixel<634) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=634 && yPixel<636) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=636 && yPixel<637) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=637 && yPixel<638) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=423 && xPixel<424 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=0 && yPixel<11) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=11 && yPixel<12) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=12 && yPixel<131) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=131 && yPixel<132) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=132 && yPixel<138) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=138 && yPixel<140) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=140 && yPixel<141) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=141 && yPixel<142) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=142 && yPixel<143) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=143 && yPixel<144) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=144 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=151 && yPixel<158) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=158 && yPixel<160) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=160 && yPixel<167) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=167 && yPixel<169) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=169 && yPixel<176) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=176 && yPixel<184) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=184 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=198 && yPixel<199) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=199 && yPixel<203) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=203 && yPixel<205) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=205 && yPixel<206) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=206 && yPixel<217) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=217 && yPixel<309) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=309 && yPixel<312) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=312 && yPixel<317) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=317 && yPixel<323) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=323 && yPixel<331) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=331 && yPixel<332) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=332 && yPixel<344) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=344 && yPixel<353) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=353 && yPixel<369) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=369 && yPixel<377) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=377 && yPixel<378) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=378 && yPixel<380) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=380 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=395 && yPixel<396) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=396 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=397 && yPixel<401) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=401 && yPixel<407) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=407 && yPixel<416) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=416 && yPixel<418) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=418 && yPixel<425) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=425 && yPixel<427) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=427 && yPixel<428) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=428 && yPixel<538) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=538 && yPixel<547) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=547 && yPixel<548) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=548 && yPixel<549) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=549 && yPixel<550) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=550 && yPixel<551) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=551 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=572 && yPixel<588) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=588 && yPixel<596) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=596 && yPixel<600) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=600 && yPixel<623) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=623 && yPixel<635) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=635 && yPixel<638) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=424 && xPixel<425 && yPixel>=638 && yPixel<639) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=0 && yPixel<12) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=12 && yPixel<63) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=63 && yPixel<64) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=64 && yPixel<141) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=141 && yPixel<146) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=146 && yPixel<151) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=151 && yPixel<154) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=154 && yPixel<197) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=197 && yPixel<198) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=198 && yPixel<200) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=200 && yPixel<203) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=203 && yPixel<206) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=206 && yPixel<334) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=334 && yPixel<336) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=336 && yPixel<339) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=339 && yPixel<345) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=345 && yPixel<354) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=354 && yPixel<369) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=369 && yPixel<377) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=377 && yPixel<379) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=379 && yPixel<381) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=381 && yPixel<393) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b10000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=393 && yPixel<395) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=395 && yPixel<397) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=397 && yPixel<399) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=399 && yPixel<405) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=405 && yPixel<423) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=423 && yPixel<429) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=429 && yPixel<431) {VGAr,VGAg,VRAb}={8'b00000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=431 && yPixel<441) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=441 && yPixel<449) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=449 && yPixel<547) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=547 && yPixel<553) {VGAr,VGAg,VRAb}={8'b10000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=553 && yPixel<554) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=554 && yPixel<556) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=556 && yPixel<558) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=558 && yPixel<564) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=564 && yPixel<566) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=566 && yPixel<570) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=570 && yPixel<571) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=571 && yPixel<572) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=572 && yPixel<586) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=586 && yPixel<587) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=587 && yPixel<594) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=594 && yPixel<595) {VGAr,VGAg,VRAb}={8'b11000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=595 && yPixel<599) {VGAr,VGAg,VRAb}={8'b10000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=599 && yPixel<601) {VGAr,VGAg,VRAb}={8'b01000000,8'b01000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=601 && yPixel<604) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=604 && yPixel<617) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=617 && yPixel<618) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=618 && yPixel<619) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b00000000};
	if(xPixel>=425 && xPixel<426 && yPixel>=619 && yPixel<639) {VGAr,VGAg,VRAb}={8'b01000000,8'b00000000,8'b01000000};

end

endmodule
