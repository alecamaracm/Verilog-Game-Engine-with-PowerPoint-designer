module PP2VerilogDrawingController(xPixel,yPixel,VGAr,VGAg,VGAb);

input [9:0]xPixel;
input[8:0]yPixel;
output [7:0]VGAr;
output [7:0]VGAg;
output [7:0]VGAb;
reg [7:0]VGAr;
reg [7:0]VGAg;
reg [7:0]VGAb;

always @(*)
begin

	//Writing backgound color
	VGAr = 8'b11111111;
	VGAg = 8'b11111111; 
	VGAb = 8'b11111111; 

	//Drawing Solid shape "Left bar"
	if(xPixel>0 && xPixel<53 && yPixel>0 && yPixel<480)
	begin
		VGAr = 8'b01000100;
		VGAg = 8'b01110010;
		VGAb = 8'b11000100;
	end

	//Drawing Solid shape "Bottom properties"
	if(xPixel>53 && xPixel<639 && yPixel>413 && yPixel<479)
	begin
		VGAr = 8'b10101111;
		VGAg = 8'b10101011;
		VGAb = 8'b10101011;
		if(xPixel<54 || xPixel>638 || yPixel<414 || yPixel>478)    //Drawing border
		begin
			VGAr = 8'b00101111;
			VGAg = 8'b01010010;
			VGAb = 8'b10001111;
		end
	end

	//Drawing Solid shape "Random Orange box"
	if(xPixel>439 && xPixel<604 && yPixel>41 && yPixel<307)
	begin
		VGAr = 8'b11000101;
		VGAg = 8'b01011010;
		VGAb = 8'b00010001;
	end

	//Drawing Solid shape "Solid purple with transparent border"
	//   --> Allowed 50% transparent render
	if(xPixel>69 && xPixel<348 && yPixel>59 && yPixel<187)
	begin
		VGAr = 8'b01110000;
		VGAg = 8'b00110000;
		VGAb = 8'b10100000;
		if(xPixel<71 || xPixel>346 || yPixel<61 || yPixel>185)    //Drawing border
		begin
			VGAr = (8'b11111111 + VGAr) / 2;
			VGAg = (8'b11011001 + VGAg) / 2;
			VGAb = (8'b01100110 + VGAb) / 2;
		end
	end

	//Drawing Solid shape "Basic transparency"
	//   --> Allowed 50% transparent render
	if(xPixel>130 && xPixel<550 && yPixel>227 && yPixel<295)
	begin
		VGAr = 8'b01010100;
		VGAg = 8'b10000010;
		VGAb = 8'b00110101;
	end

	//Drawing Solid shape "High transparency"
	//   --> Allowed 50% transparent render
	if(xPixel>369 && xPixel<470 && yPixel>130 && yPixel<198)
	begin
		VGAr = (8'b01000000 + VGAr) / 2;
		VGAg = (8'b01000000 + VGAg) / 2;
		VGAb = (8'b01000000 + VGAb) / 2;
	end

	//Drawing Solid shape "Low transparency"
	//   --> Allowed 50% transparent render
	if(xPixel>369 && xPixel<470 && yPixel>25 && yPixel<93)
	begin
		VGAr = (8'b01010100 + VGAr) / 2;
		VGAg = (8'b10000010 + VGAg) / 2;
		VGAb = (8'b00110101 + VGAb) / 2;
	end

	//Drawing picture with compression rate: 2:1
	if(yPixel>=270 && yPixel<272 && xPixel>=69 && xPixel<107) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=107 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=109 && xPixel<113) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=113 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=145 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=157 && xPixel<163) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=165 && xPixel<171) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=171 && xPixel<189) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=191 && xPixel<217) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=217 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=223 && xPixel<249) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=249 && xPixel<251) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=253 && xPixel<257) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=270 && yPixel<272 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=69 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=145 && xPixel<173) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=173 && xPixel<177) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=177 && xPixel<183) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=183 && xPixel<185) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=185 && xPixel<215) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=215 && xPixel<219) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=219 && xPixel<233) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=233 && xPixel<247) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=247 && xPixel<251) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=272 && yPixel<274 && xPixel>=253 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=69 && xPixel<127) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=131 && xPixel<143) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=143 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=161 && xPixel<175) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=175 && xPixel<187) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=187 && xPixel<193) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=193 && xPixel<215) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=215 && xPixel<217) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=217 && xPixel<223) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=223 && xPixel<227) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=227 && xPixel<249) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=274 && yPixel<276 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=69 && xPixel<125) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=125 && xPixel<127) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=127 && xPixel<129) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=129 && xPixel<141) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=141 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=155 && xPixel<159) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=163 && xPixel<175) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=175 && xPixel<185) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=185 && xPixel<199) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=199 && xPixel<203) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=203 && xPixel<207) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=207 && xPixel<215) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=215 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=223 && xPixel<241) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=276 && yPixel<278 && xPixel>=241 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=69 && xPixel<139) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=139 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=157 && xPixel<169) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=169 && xPixel<171) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=171 && xPixel<185) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=191 && xPixel<197) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=197 && xPixel<201) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=203 && xPixel<209) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=209 && xPixel<213) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=213 && xPixel<229) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=229 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=233 && xPixel<247) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=278 && yPixel<280 && xPixel>=247 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=69 && xPixel<137) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=137 && xPixel<169) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=169 && xPixel<171) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=171 && xPixel<181) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=183 && xPixel<189) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=280 && yPixel<282 && xPixel>=189 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=69 && xPixel<135) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=135 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=145 && xPixel<149) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=149 && xPixel<173) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=173 && xPixel<175) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=177 && xPixel<187) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=187 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=191 && xPixel<201) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=201 && xPixel<205) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=205 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=233 && xPixel<241) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=241 && xPixel<255) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=282 && yPixel<284 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=69 && xPixel<135) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=135 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=145 && xPixel<153) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=153 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=155 && xPixel<169) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=169 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=181 && xPixel<185) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=185 && xPixel<189) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=191 && xPixel<235) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=235 && xPixel<241) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=241 && xPixel<249) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=284 && yPixel<286 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=69 && xPixel<135) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=135 && xPixel<143) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=143 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=155 && xPixel<169) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=169 && xPixel<187) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=187 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=193 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=223 && xPixel<225) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=225 && xPixel<235) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=239 && xPixel<243) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=243 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=247 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=286 && yPixel<288 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=71 && xPixel<75) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=75 && xPixel<83) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=83 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=85 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=87 && xPixel<147) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=149 && xPixel<163) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=165 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=177 && xPixel<185) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=187 && xPixel<191) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=191 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=203 && xPixel<237) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=288 && yPixel<290 && xPixel>=241 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=69 && xPixel<75) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=75 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=81 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=87 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=157 && xPixel<163) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=163 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=177 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=191 && xPixel<195) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=195 && xPixel<197) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=197 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=203 && xPixel<209) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=209 && xPixel<239) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=290 && yPixel<292 && xPixel>=241 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=71 && xPixel<73) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=73 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=79 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=87 && xPixel<151) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=151 && xPixel<159) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=159 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=165 && xPixel<181) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=183 && xPixel<199) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=199 && xPixel<201) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=201 && xPixel<237) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=237 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=241 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=292 && yPixel<294 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=69 && xPixel<75) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=75 && xPixel<79) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=79 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=85 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=87 && xPixel<147) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=147 && xPixel<159) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=163 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=167 && xPixel<169) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=169 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=175 && xPixel<179) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=179 && xPixel<183) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=183 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=191 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=205 && xPixel<207) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=207 && xPixel<221) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=221 && xPixel<231) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=231 && xPixel<235) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=239 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=245 && xPixel<251) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=294 && yPixel<296 && xPixel>=251 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=69 && xPixel<97) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=97 && xPixel<141) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=141 && xPixel<161) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=165 && xPixel<169) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=169 && xPixel<171) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=171 && xPixel<179) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=179 && xPixel<183) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=183 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=191 && xPixel<201) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=203 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=207 && xPixel<217) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=217 && xPixel<219) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=219 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=225 && xPixel<231) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=231 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=243 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=245 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=296 && yPixel<298 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=69 && xPixel<83) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=83 && xPixel<85) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=85 && xPixel<97) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=97 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=103 && xPixel<143) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=143 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=145 && xPixel<165) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=165 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=167 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=181 && xPixel<185) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=185 && xPixel<193) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=193 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=195 && xPixel<197) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=197 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=205 && xPixel<207) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=207 && xPixel<229) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=229 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=231 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=233 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=243 && xPixel<245) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=298 && yPixel<300 && xPixel>=245 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=71 && xPixel<73) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=73 && xPixel<77) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=77 && xPixel<83) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=83 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=85 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=115 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=145 && xPixel<153) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=153 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=159 && xPixel<167) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=167 && xPixel<169) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=169 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=183 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b11000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b11000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=191 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b11000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=195 && xPixel<199) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=199 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=203 && xPixel<207) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=207 && xPixel<229) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=229 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=231 && xPixel<239) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=239 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=300 && yPixel<302 && xPixel>=245 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=69 && xPixel<83) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=83 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=87 && xPixel<97) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=97 && xPixel<99) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=99 && xPixel<117) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=117 && xPixel<129) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=129 && xPixel<131) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=131 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=145 && xPixel<149) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=151 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=157 && xPixel<165) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=165 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=181 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11000000,8'b11000000,8'b11111111};
	if(yPixel>=302 && yPixel<304 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b11000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b11000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=193 && xPixel<201) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=203 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=207 && xPixel<219) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=219 && xPixel<225) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=225 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=233 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=241 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=302 && yPixel<304 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=71 && xPixel<83) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=83 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=85 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=87 && xPixel<89) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=89 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=95 && xPixel<101) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=101 && xPixel<107) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=107 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=113 && xPixel<115) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=115 && xPixel<123) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=123 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=125 && xPixel<133) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=135 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=145 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=157 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=165 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=167 && xPixel<171) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=171 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b11000000,8'b11111111};
	if(yPixel>=304 && yPixel<306 && xPixel>=183 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b11000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=185 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=191 && xPixel<209) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=209 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=215 && xPixel<221) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=221 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=225 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=237 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=245 && xPixel<251) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=251 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=255 && xPixel<257) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=304 && yPixel<306 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=69 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=85 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=87 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=91 && xPixel<93) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=93 && xPixel<95) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=95 && xPixel<97) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=97 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=103 && xPixel<107) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=107 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=111 && xPixel<115) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=115 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=121 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=139 && xPixel<147) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=147 && xPixel<159) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=161 && xPixel<169) {VGAr,VGAg,VGAb}={8'b10000000,8'b10000000,8'b11000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=169 && xPixel<185) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=185 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=203 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=217 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=223 && xPixel<225) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=225 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=239 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=306 && yPixel<308 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=71 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=89 && xPixel<95) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=95 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=111 && xPixel<121) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=121 && xPixel<127) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=127 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=137 && xPixel<147) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=147 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=155 && xPixel<161) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=163 && xPixel<173) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=173 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=191 && xPixel<197) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=197 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=203 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=209 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=213 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=223 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=229 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=233 && xPixel<237) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=237 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=241 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=247 && xPixel<249) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=249 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b10000000};
	if(yPixel>=308 && yPixel<310 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=73 && xPixel<83) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=83 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=85 && xPixel<93) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=93 && xPixel<95) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=95 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=103 && xPixel<113) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=113 && xPixel<117) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=117 && xPixel<125) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=125 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=135 && xPixel<141) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=141 && xPixel<143) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=143 && xPixel<149) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=149 && xPixel<155) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=157 && xPixel<161) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=161 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=165 && xPixel<169) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=169 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=183 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=193 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=195 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=209 && xPixel<211) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=211 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=217 && xPixel<221) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=221 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=223 && xPixel<229) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=229 && xPixel<231) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=231 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=243 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=245 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=247 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=255 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b10000000};
	if(yPixel>=310 && yPixel<312 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=69 && xPixel<75) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=75 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=77 && xPixel<101) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=101 && xPixel<105) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=105 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=107 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=113 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=137 && xPixel<145) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=145 && xPixel<157) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=157 && xPixel<161) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=163 && xPixel<173) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=173 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=177 && xPixel<179) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=179 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=183 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=205 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=209 && xPixel<211) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=211 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=223 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=239 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=253 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=312 && yPixel<314 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=69 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=79 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=81 && xPixel<101) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=101 && xPixel<103) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=103 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=113 && xPixel<117) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=117 && xPixel<121) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b10000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=121 && xPixel<123) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=123 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=131 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=139 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=141 && xPixel<143) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=143 && xPixel<157) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=165 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=167 && xPixel<171) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=171 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=177 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=191 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=203 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=207 && xPixel<211) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=211 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=213 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=215 && xPixel<217) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=217 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=219 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=231 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=233 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=235 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=241 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=314 && yPixel<316 && xPixel>=253 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=69 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=79 && xPixel<85) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=85 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=87 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=89 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=107 && xPixel<109) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=111 && xPixel<115) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=115 && xPixel<119) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=119 && xPixel<121) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=121 && xPixel<125) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=125 && xPixel<129) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=129 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=137 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=151 && xPixel<157) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=157 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=165 && xPixel<171) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=171 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=173 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=189 && xPixel<199) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=199 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=209 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=225 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=227 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=233 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=237 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=245 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=316 && yPixel<318 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=69 && xPixel<83) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=83 && xPixel<87) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=87 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=89 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=91 && xPixel<105) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=105 && xPixel<119) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=119 && xPixel<123) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=123 && xPixel<125) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=125 && xPixel<129) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=129 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=151 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=163 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=167 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=169 && xPixel<171) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=171 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=189 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=193 && xPixel<197) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=197 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=225 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=233 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=243 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=245 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=318 && yPixel<320 && xPixel>=247 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=69 && xPixel<85) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=85 && xPixel<89) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=89 && xPixel<93) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=93 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=107 && xPixel<109) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b11000000,8'b10000000,8'b10000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=113 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=135 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=147 && xPixel<151) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=151 && xPixel<159) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=159 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=167 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=173 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=175 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=189 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=195 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=221 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=235 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=239 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=243 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=320 && yPixel<322 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=69 && xPixel<101) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=101 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=107 && xPixel<109) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=109 && xPixel<113) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b10000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=113 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b10000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=115 && xPixel<117) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=117 && xPixel<129) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=129 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=139 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=145 && xPixel<153) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=153 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=157 && xPixel<163) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=165 && xPixel<171) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=171 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=173 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=175 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=191 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=195 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=217 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=231 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=233 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=235 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=247 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b10000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=322 && yPixel<324 && xPixel>=253 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=69 && xPixel<99) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=99 && xPixel<101) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=101 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=119 && xPixel<123) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=123 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=141 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=147 && xPixel<151) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=151 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=153 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=157 && xPixel<163) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=165 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=169 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=189 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=195 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=209 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=225 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=227 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=231 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=243 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b10000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=247 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=324 && yPixel<326 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=69 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=97 && xPixel<99) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=99 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=115 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=119 && xPixel<127) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=127 && xPixel<133) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=137 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=141 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=149 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=153 && xPixel<155) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=157 && xPixel<161) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=165 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=187 && xPixel<197) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=197 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=213 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=217 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=223 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=227 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=229 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b10000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=241 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=326 && yPixel<328 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=71 && xPixel<75) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=75 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=81 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=87 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=97 && xPixel<99) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=99 && xPixel<103) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=103 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=113 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=121 && xPixel<125) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=125 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=131 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=153 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=159 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=205 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=217 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=221 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=227 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=231 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=249 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=328 && yPixel<330 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=71 && xPixel<79) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=79 && xPixel<83) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=83 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=89 && xPixel<97) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=97 && xPixel<99) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=99 && xPixel<101) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=101 && xPixel<103) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=103 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=107 && xPixel<109) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=109 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=113 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=121 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=135 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=143 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=145 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=149 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=153 && xPixel<155) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=159 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=167 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=213 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=330 && yPixel<332 && xPixel>=241 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=69 && xPixel<75) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=75 && xPixel<81) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=81 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=85 && xPixel<95) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=95 && xPixel<97) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=97 && xPixel<99) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=99 && xPixel<103) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=103 && xPixel<105) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=105 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=107 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=119 && xPixel<121) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=121 && xPixel<129) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=129 && xPixel<133) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=137 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=145 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=147 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=153 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=159 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=207 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=233 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=237 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b10000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=245 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=332 && yPixel<334 && xPixel>=247 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=73 && xPixel<79) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=79 && xPixel<87) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=87 && xPixel<91) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=91 && xPixel<99) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=99 && xPixel<105) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=105 && xPixel<109) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=109 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=113 && xPixel<115) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=115 && xPixel<121) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=121 && xPixel<125) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=125 && xPixel<127) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=131 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=137 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=147 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=207 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=217 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=219 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=227 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=231 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b10000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=241 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=334 && yPixel<336 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=73 && xPixel<77) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=77 && xPixel<79) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=79 && xPixel<93) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=93 && xPixel<99) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=99 && xPixel<105) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=105 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=115 && xPixel<119) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=119 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=135 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=147 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=153 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=165 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=169 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=177 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=205 && xPixel<211) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=211 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=213 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=223 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=225 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=229 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=239 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=243 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=245 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=336 && yPixel<338 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=77 && xPixel<79) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=79 && xPixel<81) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=81 && xPixel<85) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=85 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=119 && xPixel<125) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=125 && xPixel<127) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=127 && xPixel<129) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=129 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=135 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=145 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=149 && xPixel<161) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=161 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=165 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=167 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=195 && xPixel<199) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=199 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=209 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=219 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b10000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=223 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=233 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=237 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=243 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=338 && yPixel<340 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=77 && xPixel<81) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=81 && xPixel<83) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=83 && xPixel<89) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=89 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=125 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=135 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=147 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=153 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=203 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=205 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b11111111,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=207 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b10000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=213 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=229 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=245 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=253 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=340 && yPixel<342 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=69 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=81 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=85 && xPixel<89) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=89 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=127 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=141 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=145 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=153 && xPixel<155) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=155 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=157 && xPixel<159) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=161 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=183 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=185 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=189 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=193 && xPixel<199) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=199 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b11111111,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=205 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=223 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=225 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=235 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=239 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=251 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=342 && yPixel<344 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=69 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=79 && xPixel<89) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=89 && xPixel<93) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=93 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=95 && xPixel<117) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=117 && xPixel<133) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=137 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=141 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=145 && xPixel<163) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=163 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=169 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=173 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=175 && xPixel<177) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=177 && xPixel<179) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=179 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=185 && xPixel<197) {VGAr,VGAg,VGAb}={8'b11111111,8'b11111111,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=197 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=213 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=219 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=221 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=229 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=239 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=344 && yPixel<346 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=69 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=81 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=97 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=119 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=141 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=149 && xPixel<155) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=155 && xPixel<163) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=163 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=205 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=207 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=221 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=223 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=229 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=231 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=235 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=346 && yPixel<348 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=69 && xPixel<91) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=91 && xPixel<101) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=101 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=133 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=151 && xPixel<155) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=155 && xPixel<161) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=161 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=167 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=169 && xPixel<177) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=181 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=189 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=203 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=205 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=209 && xPixel<215) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=215 && xPixel<217) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=217 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=219 && xPixel<235) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=239 && xPixel<247) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=247 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=348 && yPixel<350 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=71 && xPixel<111) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=111 && xPixel<121) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=121 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=137 && xPixel<149) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=151 && xPixel<153) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=153 && xPixel<155) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=155 && xPixel<159) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=159 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=163 && xPixel<171) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=171 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=173 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=175 && xPixel<179) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=179 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=187 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=193 && xPixel<201) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=203 && xPixel<207) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=207 && xPixel<219) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=219 && xPixel<221) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=221 && xPixel<223) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=223 && xPixel<243) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=350 && yPixel<352 && xPixel>=243 && xPixel<259) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=69 && xPixel<149) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=149 && xPixel<173) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=173 && xPixel<177) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=177 && xPixel<185) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=187 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=193 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=195 && xPixel<197) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=197 && xPixel<201) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=201 && xPixel<209) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=209 && xPixel<245) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=352 && yPixel<354 && xPixel>=245 && xPixel<259) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=69 && xPixel<119) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=119 && xPixel<139) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=143 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=167 && xPixel<197) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=197 && xPixel<209) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=209 && xPixel<213) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=213 && xPixel<219) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=219 && xPixel<223) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b00000000};
	if(yPixel>=354 && yPixel<356 && xPixel>=223 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=73 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=81 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=95 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=125 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=133 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=143 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=151 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=157 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=187 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=191 && xPixel<197) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=197 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=209 && xPixel<211) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=211 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=221 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=231 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=235 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=356 && yPixel<358 && xPixel>=239 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=71 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=77 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=95 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=125 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=133 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=141 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=143 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=151 && xPixel<157) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=157 && xPixel<161) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=163 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=185 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=187 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=195 && xPixel<197) {VGAr,VGAg,VGAb}={8'b11111111,8'b11000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=197 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=225 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=227 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=229 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=235 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=241 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=358 && yPixel<360 && xPixel>=245 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=77 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=79 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=89 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=95 && xPixel<117) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=119 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=121 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=125 && xPixel<129) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=129 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=135 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=141 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=147 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=151 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=165 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=169 && xPixel<171) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=171 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=227 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=243 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=360 && yPixel<362 && xPixel>=253 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=77 && xPixel<81) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=81 && xPixel<93) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=93 && xPixel<99) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=99 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=115 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=121 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=125 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=135 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=141 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=149 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=151 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=169 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=239 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=243 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=362 && yPixel<364 && xPixel>=247 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=69 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=79 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=85 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=95 && xPixel<105) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=105 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=115 && xPixel<125) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=125 && xPixel<131) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=135 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=147 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=149 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=173 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=217 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=219 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=229 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=231 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=364 && yPixel<366 && xPixel>=249 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=69 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=79 && xPixel<85) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=85 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=89 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=95 && xPixel<107) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=107 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=111 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=135 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=143 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=145 && xPixel<149) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=149 && xPixel<181) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=181 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=366 && yPixel<368 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=69 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=79 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=91 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=97 && xPixel<109) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=111 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=137 && xPixel<143) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=147 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=151 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=193 && xPixel<201) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=203 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=215 && xPixel<219) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=219 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=245 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=247 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=249 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=368 && yPixel<370 && xPixel>=253 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=77 && xPixel<87) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=87 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=89 && xPixel<91) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=95 && xPixel<105) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=105 && xPixel<107) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=107 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=113 && xPixel<115) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=115 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=137 && xPixel<141) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=141 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=147 && xPixel<153) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=153 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=195 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=213 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=215 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=221 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=223 && xPixel<225) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=225 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=233 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=237 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=245 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=370 && yPixel<372 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=69 && xPixel<75) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=75 && xPixel<81) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=81 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=97 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=103 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=113 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=137 && xPixel<151) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=151 && xPixel<155) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=155 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=173 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=193 && xPixel<203) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=203 && xPixel<211) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=211 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=215 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=217 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=223 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=231 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=233 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=253 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=372 && yPixel<374 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=77 && xPixel<83) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=83 && xPixel<89) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=89 && xPixel<93) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=93 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=97 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=103 && xPixel<115) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=115 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=127 && xPixel<129) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=129 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=135 && xPixel<165) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=165 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=173 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=207 && xPixel<209) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=209 && xPixel<223) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=223 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=231 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=233 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=243 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=245 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=247 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=374 && yPixel<376 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=69 && xPixel<87) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=87 && xPixel<91) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=91 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=95 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=103 && xPixel<117) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=119 && xPixel<129) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=129 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=139 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=167 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=169 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=183 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=187 && xPixel<205) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=205 && xPixel<213) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=213 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=215 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=227 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=237 && xPixel<247) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=247 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=253 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=376 && yPixel<378 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=71 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=77 && xPixel<87) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=87 && xPixel<89) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=89 && xPixel<95) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=95 && xPixel<97) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=97 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=111 && xPixel<115) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=115 && xPixel<117) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=119 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=121 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=127 && xPixel<131) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=131 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=137 && xPixel<145) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=145 && xPixel<147) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=147 && xPixel<169) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=169 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=175 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=187 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=195 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=217 && xPixel<221) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=221 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=227 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=229 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=378 && yPixel<380 && xPixel>=243 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=69 && xPixel<89) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=89 && xPixel<93) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=93 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=97 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=103 && xPixel<115) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=115 && xPixel<117) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=117 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=135 && xPixel<139) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=139 && xPixel<155) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=155 && xPixel<159) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=159 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=193 && xPixel<207) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=207 && xPixel<211) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=211 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=215 && xPixel<217) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=217 && xPixel<227) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=227 && xPixel<233) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=233 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=243 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=251 && xPixel<253) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=253 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=380 && yPixel<382 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=69 && xPixel<97) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=97 && xPixel<103) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=103 && xPixel<113) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=113 && xPixel<119) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=119 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=139 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=165 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=167 && xPixel<171) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=171 && xPixel<175) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=175 && xPixel<181) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=181 && xPixel<189) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=191 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=193 && xPixel<197) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=197 && xPixel<199) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=199 && xPixel<201) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=203 && xPixel<211) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=211 && xPixel<215) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=215 && xPixel<217) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=217 && xPixel<235) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=235 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=243 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=249 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=382 && yPixel<384 && xPixel>=251 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=69 && xPixel<85) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=85 && xPixel<99) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=99 && xPixel<113) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=113 && xPixel<115) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=115 && xPixel<117) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=117 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=121 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=133 && xPixel<139) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=139 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=163 && xPixel<165) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=165 && xPixel<169) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=169 && xPixel<173) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=173 && xPixel<177) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=177 && xPixel<181) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=183 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=185 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=193 && xPixel<199) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=199 && xPixel<201) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=203 && xPixel<231) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=231 && xPixel<237) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=237 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=241 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11111111,8'b10000000,8'b01000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=243 && xPixel<249) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=249 && xPixel<251) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b01000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=251 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=384 && yPixel<386 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=73 && xPixel<75) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=75 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=81 && xPixel<83) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=83 && xPixel<87) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=87 && xPixel<99) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=99 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=113 && xPixel<115) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=115 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=127 && xPixel<129) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=129 && xPixel<131) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=133 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=137 && xPixel<143) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=143 && xPixel<147) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=147 && xPixel<151) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=151 && xPixel<165) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=165 && xPixel<167) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=167 && xPixel<181) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=181 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=183 && xPixel<193) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=193 && xPixel<199) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=199 && xPixel<201) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=201 && xPixel<203) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=203 && xPixel<209) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=209 && xPixel<211) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=211 && xPixel<245) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=245 && xPixel<255) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=255 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=386 && yPixel<388 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11111111,8'b01000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=69 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=77 && xPixel<85) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=85 && xPixel<103) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=103 && xPixel<107) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=107 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=113 && xPixel<117) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=119 && xPixel<121) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=121 && xPixel<123) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=123 && xPixel<127) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=127 && xPixel<129) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=129 && xPixel<133) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=133 && xPixel<145) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=145 && xPixel<151) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=151 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=167 && xPixel<171) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=171 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=175 && xPixel<181) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=181 && xPixel<185) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=185 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=191 && xPixel<205) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=205 && xPixel<209) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=209 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=223 && xPixel<229) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=229 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=233 && xPixel<239) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=239 && xPixel<243) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=243 && xPixel<249) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=249 && xPixel<257) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=388 && yPixel<390 && xPixel>=257 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=73 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=77 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=81 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=111 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=113 && xPixel<117) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=119 && xPixel<125) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=125 && xPixel<129) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=129 && xPixel<131) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=131 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=139 && xPixel<143) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=143 && xPixel<145) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=145 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=155 && xPixel<171) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=171 && xPixel<175) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=175 && xPixel<187) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=187 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=191 && xPixel<203) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=203 && xPixel<229) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=229 && xPixel<239) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=390 && yPixel<392 && xPixel>=239 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=69 && xPixel<71) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=71 && xPixel<77) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=77 && xPixel<81) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=81 && xPixel<111) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=111 && xPixel<115) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=115 && xPixel<117) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=119 && xPixel<121) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=121 && xPixel<123) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=123 && xPixel<125) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=125 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=137 && xPixel<139) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=139 && xPixel<141) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=141 && xPixel<163) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=163 && xPixel<167) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=167 && xPixel<171) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=171 && xPixel<173) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=173 && xPixel<183) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=183 && xPixel<187) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=187 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=195 && xPixel<205) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=205 && xPixel<211) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=211 && xPixel<213) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=213 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=223 && xPixel<243) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=243 && xPixel<247) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=247 && xPixel<249) {VGAr,VGAg,VGAb}={8'b01000000,8'b01000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=249 && xPixel<253) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=392 && yPixel<394 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=69 && xPixel<75) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=75 && xPixel<79) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=79 && xPixel<103) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=103 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=109 && xPixel<111) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=111 && xPixel<121) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=121 && xPixel<123) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=123 && xPixel<127) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=127 && xPixel<129) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=129 && xPixel<133) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=133 && xPixel<135) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=135 && xPixel<137) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=137 && xPixel<143) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=143 && xPixel<145) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=145 && xPixel<155) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=155 && xPixel<159) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=159 && xPixel<161) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=161 && xPixel<163) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=163 && xPixel<167) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=167 && xPixel<169) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=169 && xPixel<179) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=179 && xPixel<185) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=185 && xPixel<191) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=191 && xPixel<195) {VGAr,VGAg,VGAb}={8'b11000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=195 && xPixel<207) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=207 && xPixel<219) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=219 && xPixel<223) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=223 && xPixel<227) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=227 && xPixel<231) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=231 && xPixel<233) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=233 && xPixel<235) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=235 && xPixel<237) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=237 && xPixel<239) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=239 && xPixel<245) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=245 && xPixel<251) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=394 && yPixel<396 && xPixel>=251 && xPixel<259) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b01000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=69 && xPixel<73) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=73 && xPixel<109) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=109 && xPixel<113) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=113 && xPixel<117) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=117 && xPixel<119) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=119 && xPixel<123) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=123 && xPixel<131) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=131 && xPixel<153) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=153 && xPixel<161) {VGAr,VGAg,VGAb}={8'b00000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=161 && xPixel<167) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=167 && xPixel<175) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=175 && xPixel<183) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=183 && xPixel<187) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=187 && xPixel<189) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=189 && xPixel<191) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=191 && xPixel<201) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=201 && xPixel<213) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=213 && xPixel<221) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=221 && xPixel<229) {VGAr,VGAg,VGAb}={8'b10000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=229 && xPixel<231) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=231 && xPixel<241) {VGAr,VGAg,VGAb}={8'b11000000,8'b01000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=241 && xPixel<245) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=245 && xPixel<249) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=249 && xPixel<253) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b00000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=253 && xPixel<255) {VGAr,VGAg,VGAb}={8'b01000000,8'b00000000,8'b01000000};
	if(yPixel>=396 && yPixel<398 && xPixel>=255 && xPixel<259) {VGAr,VGAg,VGAb}={8'b10000000,8'b01000000,8'b01000000};

end

endmodule
